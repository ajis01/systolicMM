module EnumOps(
  input  [6:0] io_x,
  input  [6:0] io_y,
  output       io_lt,
  output       io_le,
  output       io_gt,
  output       io_ge,
  output       io_eq,
  output       io_ne
);
  assign io_lt = io_x < io_y; // @[StrongEnum.scala 98:9]
  assign io_le = io_x <= io_y; // @[StrongEnum.scala 99:9]
  assign io_gt = io_x > io_y; // @[StrongEnum.scala 100:9]
  assign io_ge = io_x >= io_y; // @[StrongEnum.scala 101:9]
  assign io_eq = io_x == io_y; // @[StrongEnum.scala 102:9]
  assign io_ne = io_x != io_y; // @[StrongEnum.scala 103:9]
endmodule
module EnumOpsTester(
  input   clock,
  input   reset
);
  wire [6:0] EnumOps_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_1_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_1_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_1_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_1_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_1_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_1_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_1_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_1_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_2_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_2_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_2_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_2_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_2_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_2_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_2_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_2_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_3_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_3_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_3_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_3_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_3_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_3_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_3_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_3_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_4_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_4_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_4_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_4_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_4_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_4_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_4_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_4_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_5_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_5_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_5_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_5_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_5_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_5_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_5_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_5_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_6_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_6_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_6_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_6_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_6_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_6_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_6_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_6_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_7_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_7_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_7_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_7_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_7_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_7_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_7_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_7_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_8_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_8_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_8_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_8_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_8_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_8_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_8_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_8_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_9_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_9_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_9_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_9_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_9_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_9_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_9_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_9_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_10_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_10_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_10_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_10_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_10_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_10_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_10_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_10_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_11_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_11_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_11_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_11_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_11_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_11_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_11_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_11_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_12_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_12_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_12_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_12_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_12_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_12_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_12_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_12_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_13_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_13_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_13_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_13_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_13_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_13_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_13_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_13_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_14_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_14_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_14_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_14_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_14_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_14_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_14_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_14_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_15_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_15_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_15_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_15_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_15_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_15_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_15_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_15_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_16_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_16_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_16_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_16_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_16_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_16_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_16_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_16_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_17_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_17_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_17_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_17_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_17_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_17_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_17_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_17_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_18_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_18_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_18_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_18_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_18_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_18_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_18_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_18_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_19_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_19_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_19_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_19_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_19_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_19_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_19_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_19_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_20_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_20_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_20_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_20_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_20_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_20_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_20_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_20_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_21_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_21_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_21_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_21_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_21_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_21_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_21_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_21_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_22_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_22_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_22_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_22_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_22_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_22_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_22_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_22_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_23_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_23_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_23_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_23_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_23_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_23_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_23_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_23_io_ne; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_24_io_x; // @[StrongEnum.scala 199:21]
  wire [6:0] EnumOps_24_io_y; // @[StrongEnum.scala 199:21]
  wire  EnumOps_24_io_lt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_24_io_le; // @[StrongEnum.scala 199:21]
  wire  EnumOps_24_io_gt; // @[StrongEnum.scala 199:21]
  wire  EnumOps_24_io_ge; // @[StrongEnum.scala 199:21]
  wire  EnumOps_24_io_eq; // @[StrongEnum.scala 199:21]
  wire  EnumOps_24_io_ne; // @[StrongEnum.scala 199:21]
  wire  _T_3; // @[StrongEnum.scala 203:22]
  wire  _T_5; // @[StrongEnum.scala 203:11]
  wire  _T_6; // @[StrongEnum.scala 203:11]
  wire  _T_10; // @[StrongEnum.scala 204:22]
  wire  _T_12; // @[StrongEnum.scala 204:11]
  wire  _T_13; // @[StrongEnum.scala 204:11]
  wire  _T_17; // @[StrongEnum.scala 205:22]
  wire  _T_19; // @[StrongEnum.scala 205:11]
  wire  _T_20; // @[StrongEnum.scala 205:11]
  wire  _T_24; // @[StrongEnum.scala 206:22]
  wire  _T_26; // @[StrongEnum.scala 206:11]
  wire  _T_27; // @[StrongEnum.scala 206:11]
  wire  _T_31; // @[StrongEnum.scala 207:22]
  wire  _T_33; // @[StrongEnum.scala 207:11]
  wire  _T_34; // @[StrongEnum.scala 207:11]
  wire  _T_38; // @[StrongEnum.scala 208:22]
  wire  _T_40; // @[StrongEnum.scala 208:11]
  wire  _T_41; // @[StrongEnum.scala 208:11]
  wire  _T_45; // @[StrongEnum.scala 203:22]
  wire  _T_47; // @[StrongEnum.scala 203:11]
  wire  _T_48; // @[StrongEnum.scala 203:11]
  wire  _T_52; // @[StrongEnum.scala 204:22]
  wire  _T_54; // @[StrongEnum.scala 204:11]
  wire  _T_55; // @[StrongEnum.scala 204:11]
  wire  _T_59; // @[StrongEnum.scala 205:22]
  wire  _T_61; // @[StrongEnum.scala 205:11]
  wire  _T_62; // @[StrongEnum.scala 205:11]
  wire  _T_66; // @[StrongEnum.scala 206:22]
  wire  _T_68; // @[StrongEnum.scala 206:11]
  wire  _T_69; // @[StrongEnum.scala 206:11]
  wire  _T_73; // @[StrongEnum.scala 207:22]
  wire  _T_75; // @[StrongEnum.scala 207:11]
  wire  _T_76; // @[StrongEnum.scala 207:11]
  wire  _T_80; // @[StrongEnum.scala 208:22]
  wire  _T_82; // @[StrongEnum.scala 208:11]
  wire  _T_83; // @[StrongEnum.scala 208:11]
  wire  _T_87; // @[StrongEnum.scala 203:22]
  wire  _T_89; // @[StrongEnum.scala 203:11]
  wire  _T_90; // @[StrongEnum.scala 203:11]
  wire  _T_94; // @[StrongEnum.scala 204:22]
  wire  _T_96; // @[StrongEnum.scala 204:11]
  wire  _T_97; // @[StrongEnum.scala 204:11]
  wire  _T_101; // @[StrongEnum.scala 205:22]
  wire  _T_103; // @[StrongEnum.scala 205:11]
  wire  _T_104; // @[StrongEnum.scala 205:11]
  wire  _T_108; // @[StrongEnum.scala 206:22]
  wire  _T_110; // @[StrongEnum.scala 206:11]
  wire  _T_111; // @[StrongEnum.scala 206:11]
  wire  _T_115; // @[StrongEnum.scala 207:22]
  wire  _T_117; // @[StrongEnum.scala 207:11]
  wire  _T_118; // @[StrongEnum.scala 207:11]
  wire  _T_122; // @[StrongEnum.scala 208:22]
  wire  _T_124; // @[StrongEnum.scala 208:11]
  wire  _T_125; // @[StrongEnum.scala 208:11]
  wire  _T_129; // @[StrongEnum.scala 203:22]
  wire  _T_131; // @[StrongEnum.scala 203:11]
  wire  _T_132; // @[StrongEnum.scala 203:11]
  wire  _T_136; // @[StrongEnum.scala 204:22]
  wire  _T_138; // @[StrongEnum.scala 204:11]
  wire  _T_139; // @[StrongEnum.scala 204:11]
  wire  _T_143; // @[StrongEnum.scala 205:22]
  wire  _T_145; // @[StrongEnum.scala 205:11]
  wire  _T_146; // @[StrongEnum.scala 205:11]
  wire  _T_150; // @[StrongEnum.scala 206:22]
  wire  _T_152; // @[StrongEnum.scala 206:11]
  wire  _T_153; // @[StrongEnum.scala 206:11]
  wire  _T_157; // @[StrongEnum.scala 207:22]
  wire  _T_159; // @[StrongEnum.scala 207:11]
  wire  _T_160; // @[StrongEnum.scala 207:11]
  wire  _T_164; // @[StrongEnum.scala 208:22]
  wire  _T_166; // @[StrongEnum.scala 208:11]
  wire  _T_167; // @[StrongEnum.scala 208:11]
  wire  _T_171; // @[StrongEnum.scala 203:22]
  wire  _T_173; // @[StrongEnum.scala 203:11]
  wire  _T_174; // @[StrongEnum.scala 203:11]
  wire  _T_178; // @[StrongEnum.scala 204:22]
  wire  _T_180; // @[StrongEnum.scala 204:11]
  wire  _T_181; // @[StrongEnum.scala 204:11]
  wire  _T_185; // @[StrongEnum.scala 205:22]
  wire  _T_187; // @[StrongEnum.scala 205:11]
  wire  _T_188; // @[StrongEnum.scala 205:11]
  wire  _T_192; // @[StrongEnum.scala 206:22]
  wire  _T_194; // @[StrongEnum.scala 206:11]
  wire  _T_195; // @[StrongEnum.scala 206:11]
  wire  _T_199; // @[StrongEnum.scala 207:22]
  wire  _T_201; // @[StrongEnum.scala 207:11]
  wire  _T_202; // @[StrongEnum.scala 207:11]
  wire  _T_206; // @[StrongEnum.scala 208:22]
  wire  _T_208; // @[StrongEnum.scala 208:11]
  wire  _T_209; // @[StrongEnum.scala 208:11]
  wire  _T_213; // @[StrongEnum.scala 203:22]
  wire  _T_215; // @[StrongEnum.scala 203:11]
  wire  _T_216; // @[StrongEnum.scala 203:11]
  wire  _T_220; // @[StrongEnum.scala 204:22]
  wire  _T_222; // @[StrongEnum.scala 204:11]
  wire  _T_223; // @[StrongEnum.scala 204:11]
  wire  _T_227; // @[StrongEnum.scala 205:22]
  wire  _T_229; // @[StrongEnum.scala 205:11]
  wire  _T_230; // @[StrongEnum.scala 205:11]
  wire  _T_234; // @[StrongEnum.scala 206:22]
  wire  _T_236; // @[StrongEnum.scala 206:11]
  wire  _T_237; // @[StrongEnum.scala 206:11]
  wire  _T_241; // @[StrongEnum.scala 207:22]
  wire  _T_243; // @[StrongEnum.scala 207:11]
  wire  _T_244; // @[StrongEnum.scala 207:11]
  wire  _T_248; // @[StrongEnum.scala 208:22]
  wire  _T_250; // @[StrongEnum.scala 208:11]
  wire  _T_251; // @[StrongEnum.scala 208:11]
  wire  _T_255; // @[StrongEnum.scala 203:22]
  wire  _T_257; // @[StrongEnum.scala 203:11]
  wire  _T_258; // @[StrongEnum.scala 203:11]
  wire  _T_262; // @[StrongEnum.scala 204:22]
  wire  _T_264; // @[StrongEnum.scala 204:11]
  wire  _T_265; // @[StrongEnum.scala 204:11]
  wire  _T_269; // @[StrongEnum.scala 205:22]
  wire  _T_271; // @[StrongEnum.scala 205:11]
  wire  _T_272; // @[StrongEnum.scala 205:11]
  wire  _T_276; // @[StrongEnum.scala 206:22]
  wire  _T_278; // @[StrongEnum.scala 206:11]
  wire  _T_279; // @[StrongEnum.scala 206:11]
  wire  _T_283; // @[StrongEnum.scala 207:22]
  wire  _T_285; // @[StrongEnum.scala 207:11]
  wire  _T_286; // @[StrongEnum.scala 207:11]
  wire  _T_290; // @[StrongEnum.scala 208:22]
  wire  _T_292; // @[StrongEnum.scala 208:11]
  wire  _T_293; // @[StrongEnum.scala 208:11]
  wire  _T_297; // @[StrongEnum.scala 203:22]
  wire  _T_299; // @[StrongEnum.scala 203:11]
  wire  _T_300; // @[StrongEnum.scala 203:11]
  wire  _T_304; // @[StrongEnum.scala 204:22]
  wire  _T_306; // @[StrongEnum.scala 204:11]
  wire  _T_307; // @[StrongEnum.scala 204:11]
  wire  _T_311; // @[StrongEnum.scala 205:22]
  wire  _T_313; // @[StrongEnum.scala 205:11]
  wire  _T_314; // @[StrongEnum.scala 205:11]
  wire  _T_318; // @[StrongEnum.scala 206:22]
  wire  _T_320; // @[StrongEnum.scala 206:11]
  wire  _T_321; // @[StrongEnum.scala 206:11]
  wire  _T_325; // @[StrongEnum.scala 207:22]
  wire  _T_327; // @[StrongEnum.scala 207:11]
  wire  _T_328; // @[StrongEnum.scala 207:11]
  wire  _T_332; // @[StrongEnum.scala 208:22]
  wire  _T_334; // @[StrongEnum.scala 208:11]
  wire  _T_335; // @[StrongEnum.scala 208:11]
  wire  _T_339; // @[StrongEnum.scala 203:22]
  wire  _T_341; // @[StrongEnum.scala 203:11]
  wire  _T_342; // @[StrongEnum.scala 203:11]
  wire  _T_346; // @[StrongEnum.scala 204:22]
  wire  _T_348; // @[StrongEnum.scala 204:11]
  wire  _T_349; // @[StrongEnum.scala 204:11]
  wire  _T_353; // @[StrongEnum.scala 205:22]
  wire  _T_355; // @[StrongEnum.scala 205:11]
  wire  _T_356; // @[StrongEnum.scala 205:11]
  wire  _T_360; // @[StrongEnum.scala 206:22]
  wire  _T_362; // @[StrongEnum.scala 206:11]
  wire  _T_363; // @[StrongEnum.scala 206:11]
  wire  _T_367; // @[StrongEnum.scala 207:22]
  wire  _T_369; // @[StrongEnum.scala 207:11]
  wire  _T_370; // @[StrongEnum.scala 207:11]
  wire  _T_374; // @[StrongEnum.scala 208:22]
  wire  _T_376; // @[StrongEnum.scala 208:11]
  wire  _T_377; // @[StrongEnum.scala 208:11]
  wire  _T_381; // @[StrongEnum.scala 203:22]
  wire  _T_383; // @[StrongEnum.scala 203:11]
  wire  _T_384; // @[StrongEnum.scala 203:11]
  wire  _T_388; // @[StrongEnum.scala 204:22]
  wire  _T_390; // @[StrongEnum.scala 204:11]
  wire  _T_391; // @[StrongEnum.scala 204:11]
  wire  _T_395; // @[StrongEnum.scala 205:22]
  wire  _T_397; // @[StrongEnum.scala 205:11]
  wire  _T_398; // @[StrongEnum.scala 205:11]
  wire  _T_402; // @[StrongEnum.scala 206:22]
  wire  _T_404; // @[StrongEnum.scala 206:11]
  wire  _T_405; // @[StrongEnum.scala 206:11]
  wire  _T_409; // @[StrongEnum.scala 207:22]
  wire  _T_411; // @[StrongEnum.scala 207:11]
  wire  _T_412; // @[StrongEnum.scala 207:11]
  wire  _T_416; // @[StrongEnum.scala 208:22]
  wire  _T_418; // @[StrongEnum.scala 208:11]
  wire  _T_419; // @[StrongEnum.scala 208:11]
  wire  _T_423; // @[StrongEnum.scala 203:22]
  wire  _T_425; // @[StrongEnum.scala 203:11]
  wire  _T_426; // @[StrongEnum.scala 203:11]
  wire  _T_430; // @[StrongEnum.scala 204:22]
  wire  _T_432; // @[StrongEnum.scala 204:11]
  wire  _T_433; // @[StrongEnum.scala 204:11]
  wire  _T_437; // @[StrongEnum.scala 205:22]
  wire  _T_439; // @[StrongEnum.scala 205:11]
  wire  _T_440; // @[StrongEnum.scala 205:11]
  wire  _T_444; // @[StrongEnum.scala 206:22]
  wire  _T_446; // @[StrongEnum.scala 206:11]
  wire  _T_447; // @[StrongEnum.scala 206:11]
  wire  _T_451; // @[StrongEnum.scala 207:22]
  wire  _T_453; // @[StrongEnum.scala 207:11]
  wire  _T_454; // @[StrongEnum.scala 207:11]
  wire  _T_458; // @[StrongEnum.scala 208:22]
  wire  _T_460; // @[StrongEnum.scala 208:11]
  wire  _T_461; // @[StrongEnum.scala 208:11]
  wire  _T_465; // @[StrongEnum.scala 203:22]
  wire  _T_467; // @[StrongEnum.scala 203:11]
  wire  _T_468; // @[StrongEnum.scala 203:11]
  wire  _T_472; // @[StrongEnum.scala 204:22]
  wire  _T_474; // @[StrongEnum.scala 204:11]
  wire  _T_475; // @[StrongEnum.scala 204:11]
  wire  _T_479; // @[StrongEnum.scala 205:22]
  wire  _T_481; // @[StrongEnum.scala 205:11]
  wire  _T_482; // @[StrongEnum.scala 205:11]
  wire  _T_486; // @[StrongEnum.scala 206:22]
  wire  _T_488; // @[StrongEnum.scala 206:11]
  wire  _T_489; // @[StrongEnum.scala 206:11]
  wire  _T_493; // @[StrongEnum.scala 207:22]
  wire  _T_495; // @[StrongEnum.scala 207:11]
  wire  _T_496; // @[StrongEnum.scala 207:11]
  wire  _T_500; // @[StrongEnum.scala 208:22]
  wire  _T_502; // @[StrongEnum.scala 208:11]
  wire  _T_503; // @[StrongEnum.scala 208:11]
  wire  _T_507; // @[StrongEnum.scala 203:22]
  wire  _T_509; // @[StrongEnum.scala 203:11]
  wire  _T_510; // @[StrongEnum.scala 203:11]
  wire  _T_514; // @[StrongEnum.scala 204:22]
  wire  _T_516; // @[StrongEnum.scala 204:11]
  wire  _T_517; // @[StrongEnum.scala 204:11]
  wire  _T_521; // @[StrongEnum.scala 205:22]
  wire  _T_523; // @[StrongEnum.scala 205:11]
  wire  _T_524; // @[StrongEnum.scala 205:11]
  wire  _T_528; // @[StrongEnum.scala 206:22]
  wire  _T_530; // @[StrongEnum.scala 206:11]
  wire  _T_531; // @[StrongEnum.scala 206:11]
  wire  _T_535; // @[StrongEnum.scala 207:22]
  wire  _T_537; // @[StrongEnum.scala 207:11]
  wire  _T_538; // @[StrongEnum.scala 207:11]
  wire  _T_542; // @[StrongEnum.scala 208:22]
  wire  _T_544; // @[StrongEnum.scala 208:11]
  wire  _T_545; // @[StrongEnum.scala 208:11]
  wire  _T_549; // @[StrongEnum.scala 203:22]
  wire  _T_551; // @[StrongEnum.scala 203:11]
  wire  _T_552; // @[StrongEnum.scala 203:11]
  wire  _T_556; // @[StrongEnum.scala 204:22]
  wire  _T_558; // @[StrongEnum.scala 204:11]
  wire  _T_559; // @[StrongEnum.scala 204:11]
  wire  _T_563; // @[StrongEnum.scala 205:22]
  wire  _T_565; // @[StrongEnum.scala 205:11]
  wire  _T_566; // @[StrongEnum.scala 205:11]
  wire  _T_570; // @[StrongEnum.scala 206:22]
  wire  _T_572; // @[StrongEnum.scala 206:11]
  wire  _T_573; // @[StrongEnum.scala 206:11]
  wire  _T_577; // @[StrongEnum.scala 207:22]
  wire  _T_579; // @[StrongEnum.scala 207:11]
  wire  _T_580; // @[StrongEnum.scala 207:11]
  wire  _T_584; // @[StrongEnum.scala 208:22]
  wire  _T_586; // @[StrongEnum.scala 208:11]
  wire  _T_587; // @[StrongEnum.scala 208:11]
  wire  _T_591; // @[StrongEnum.scala 203:22]
  wire  _T_593; // @[StrongEnum.scala 203:11]
  wire  _T_594; // @[StrongEnum.scala 203:11]
  wire  _T_598; // @[StrongEnum.scala 204:22]
  wire  _T_600; // @[StrongEnum.scala 204:11]
  wire  _T_601; // @[StrongEnum.scala 204:11]
  wire  _T_605; // @[StrongEnum.scala 205:22]
  wire  _T_607; // @[StrongEnum.scala 205:11]
  wire  _T_608; // @[StrongEnum.scala 205:11]
  wire  _T_612; // @[StrongEnum.scala 206:22]
  wire  _T_614; // @[StrongEnum.scala 206:11]
  wire  _T_615; // @[StrongEnum.scala 206:11]
  wire  _T_619; // @[StrongEnum.scala 207:22]
  wire  _T_621; // @[StrongEnum.scala 207:11]
  wire  _T_622; // @[StrongEnum.scala 207:11]
  wire  _T_626; // @[StrongEnum.scala 208:22]
  wire  _T_628; // @[StrongEnum.scala 208:11]
  wire  _T_629; // @[StrongEnum.scala 208:11]
  wire  _T_633; // @[StrongEnum.scala 203:22]
  wire  _T_635; // @[StrongEnum.scala 203:11]
  wire  _T_636; // @[StrongEnum.scala 203:11]
  wire  _T_640; // @[StrongEnum.scala 204:22]
  wire  _T_642; // @[StrongEnum.scala 204:11]
  wire  _T_643; // @[StrongEnum.scala 204:11]
  wire  _T_647; // @[StrongEnum.scala 205:22]
  wire  _T_649; // @[StrongEnum.scala 205:11]
  wire  _T_650; // @[StrongEnum.scala 205:11]
  wire  _T_654; // @[StrongEnum.scala 206:22]
  wire  _T_656; // @[StrongEnum.scala 206:11]
  wire  _T_657; // @[StrongEnum.scala 206:11]
  wire  _T_661; // @[StrongEnum.scala 207:22]
  wire  _T_663; // @[StrongEnum.scala 207:11]
  wire  _T_664; // @[StrongEnum.scala 207:11]
  wire  _T_668; // @[StrongEnum.scala 208:22]
  wire  _T_670; // @[StrongEnum.scala 208:11]
  wire  _T_671; // @[StrongEnum.scala 208:11]
  wire  _T_675; // @[StrongEnum.scala 203:22]
  wire  _T_677; // @[StrongEnum.scala 203:11]
  wire  _T_678; // @[StrongEnum.scala 203:11]
  wire  _T_682; // @[StrongEnum.scala 204:22]
  wire  _T_684; // @[StrongEnum.scala 204:11]
  wire  _T_685; // @[StrongEnum.scala 204:11]
  wire  _T_689; // @[StrongEnum.scala 205:22]
  wire  _T_691; // @[StrongEnum.scala 205:11]
  wire  _T_692; // @[StrongEnum.scala 205:11]
  wire  _T_696; // @[StrongEnum.scala 206:22]
  wire  _T_698; // @[StrongEnum.scala 206:11]
  wire  _T_699; // @[StrongEnum.scala 206:11]
  wire  _T_703; // @[StrongEnum.scala 207:22]
  wire  _T_705; // @[StrongEnum.scala 207:11]
  wire  _T_706; // @[StrongEnum.scala 207:11]
  wire  _T_710; // @[StrongEnum.scala 208:22]
  wire  _T_712; // @[StrongEnum.scala 208:11]
  wire  _T_713; // @[StrongEnum.scala 208:11]
  wire  _T_717; // @[StrongEnum.scala 203:22]
  wire  _T_719; // @[StrongEnum.scala 203:11]
  wire  _T_720; // @[StrongEnum.scala 203:11]
  wire  _T_724; // @[StrongEnum.scala 204:22]
  wire  _T_726; // @[StrongEnum.scala 204:11]
  wire  _T_727; // @[StrongEnum.scala 204:11]
  wire  _T_731; // @[StrongEnum.scala 205:22]
  wire  _T_733; // @[StrongEnum.scala 205:11]
  wire  _T_734; // @[StrongEnum.scala 205:11]
  wire  _T_738; // @[StrongEnum.scala 206:22]
  wire  _T_740; // @[StrongEnum.scala 206:11]
  wire  _T_741; // @[StrongEnum.scala 206:11]
  wire  _T_745; // @[StrongEnum.scala 207:22]
  wire  _T_747; // @[StrongEnum.scala 207:11]
  wire  _T_748; // @[StrongEnum.scala 207:11]
  wire  _T_752; // @[StrongEnum.scala 208:22]
  wire  _T_754; // @[StrongEnum.scala 208:11]
  wire  _T_755; // @[StrongEnum.scala 208:11]
  wire  _T_759; // @[StrongEnum.scala 203:22]
  wire  _T_761; // @[StrongEnum.scala 203:11]
  wire  _T_762; // @[StrongEnum.scala 203:11]
  wire  _T_766; // @[StrongEnum.scala 204:22]
  wire  _T_768; // @[StrongEnum.scala 204:11]
  wire  _T_769; // @[StrongEnum.scala 204:11]
  wire  _T_773; // @[StrongEnum.scala 205:22]
  wire  _T_775; // @[StrongEnum.scala 205:11]
  wire  _T_776; // @[StrongEnum.scala 205:11]
  wire  _T_780; // @[StrongEnum.scala 206:22]
  wire  _T_782; // @[StrongEnum.scala 206:11]
  wire  _T_783; // @[StrongEnum.scala 206:11]
  wire  _T_787; // @[StrongEnum.scala 207:22]
  wire  _T_789; // @[StrongEnum.scala 207:11]
  wire  _T_790; // @[StrongEnum.scala 207:11]
  wire  _T_794; // @[StrongEnum.scala 208:22]
  wire  _T_796; // @[StrongEnum.scala 208:11]
  wire  _T_797; // @[StrongEnum.scala 208:11]
  wire  _T_801; // @[StrongEnum.scala 203:22]
  wire  _T_803; // @[StrongEnum.scala 203:11]
  wire  _T_804; // @[StrongEnum.scala 203:11]
  wire  _T_808; // @[StrongEnum.scala 204:22]
  wire  _T_810; // @[StrongEnum.scala 204:11]
  wire  _T_811; // @[StrongEnum.scala 204:11]
  wire  _T_815; // @[StrongEnum.scala 205:22]
  wire  _T_817; // @[StrongEnum.scala 205:11]
  wire  _T_818; // @[StrongEnum.scala 205:11]
  wire  _T_822; // @[StrongEnum.scala 206:22]
  wire  _T_824; // @[StrongEnum.scala 206:11]
  wire  _T_825; // @[StrongEnum.scala 206:11]
  wire  _T_829; // @[StrongEnum.scala 207:22]
  wire  _T_831; // @[StrongEnum.scala 207:11]
  wire  _T_832; // @[StrongEnum.scala 207:11]
  wire  _T_836; // @[StrongEnum.scala 208:22]
  wire  _T_838; // @[StrongEnum.scala 208:11]
  wire  _T_839; // @[StrongEnum.scala 208:11]
  wire  _T_843; // @[StrongEnum.scala 203:22]
  wire  _T_845; // @[StrongEnum.scala 203:11]
  wire  _T_846; // @[StrongEnum.scala 203:11]
  wire  _T_850; // @[StrongEnum.scala 204:22]
  wire  _T_852; // @[StrongEnum.scala 204:11]
  wire  _T_853; // @[StrongEnum.scala 204:11]
  wire  _T_857; // @[StrongEnum.scala 205:22]
  wire  _T_859; // @[StrongEnum.scala 205:11]
  wire  _T_860; // @[StrongEnum.scala 205:11]
  wire  _T_864; // @[StrongEnum.scala 206:22]
  wire  _T_866; // @[StrongEnum.scala 206:11]
  wire  _T_867; // @[StrongEnum.scala 206:11]
  wire  _T_871; // @[StrongEnum.scala 207:22]
  wire  _T_873; // @[StrongEnum.scala 207:11]
  wire  _T_874; // @[StrongEnum.scala 207:11]
  wire  _T_878; // @[StrongEnum.scala 208:22]
  wire  _T_880; // @[StrongEnum.scala 208:11]
  wire  _T_881; // @[StrongEnum.scala 208:11]
  wire  _T_885; // @[StrongEnum.scala 203:22]
  wire  _T_887; // @[StrongEnum.scala 203:11]
  wire  _T_888; // @[StrongEnum.scala 203:11]
  wire  _T_892; // @[StrongEnum.scala 204:22]
  wire  _T_894; // @[StrongEnum.scala 204:11]
  wire  _T_895; // @[StrongEnum.scala 204:11]
  wire  _T_899; // @[StrongEnum.scala 205:22]
  wire  _T_901; // @[StrongEnum.scala 205:11]
  wire  _T_902; // @[StrongEnum.scala 205:11]
  wire  _T_906; // @[StrongEnum.scala 206:22]
  wire  _T_908; // @[StrongEnum.scala 206:11]
  wire  _T_909; // @[StrongEnum.scala 206:11]
  wire  _T_913; // @[StrongEnum.scala 207:22]
  wire  _T_915; // @[StrongEnum.scala 207:11]
  wire  _T_916; // @[StrongEnum.scala 207:11]
  wire  _T_920; // @[StrongEnum.scala 208:22]
  wire  _T_922; // @[StrongEnum.scala 208:11]
  wire  _T_923; // @[StrongEnum.scala 208:11]
  wire  _T_927; // @[StrongEnum.scala 203:22]
  wire  _T_929; // @[StrongEnum.scala 203:11]
  wire  _T_930; // @[StrongEnum.scala 203:11]
  wire  _T_934; // @[StrongEnum.scala 204:22]
  wire  _T_936; // @[StrongEnum.scala 204:11]
  wire  _T_937; // @[StrongEnum.scala 204:11]
  wire  _T_941; // @[StrongEnum.scala 205:22]
  wire  _T_943; // @[StrongEnum.scala 205:11]
  wire  _T_944; // @[StrongEnum.scala 205:11]
  wire  _T_948; // @[StrongEnum.scala 206:22]
  wire  _T_950; // @[StrongEnum.scala 206:11]
  wire  _T_951; // @[StrongEnum.scala 206:11]
  wire  _T_955; // @[StrongEnum.scala 207:22]
  wire  _T_957; // @[StrongEnum.scala 207:11]
  wire  _T_958; // @[StrongEnum.scala 207:11]
  wire  _T_962; // @[StrongEnum.scala 208:22]
  wire  _T_964; // @[StrongEnum.scala 208:11]
  wire  _T_965; // @[StrongEnum.scala 208:11]
  wire  _T_969; // @[StrongEnum.scala 203:22]
  wire  _T_971; // @[StrongEnum.scala 203:11]
  wire  _T_972; // @[StrongEnum.scala 203:11]
  wire  _T_976; // @[StrongEnum.scala 204:22]
  wire  _T_978; // @[StrongEnum.scala 204:11]
  wire  _T_979; // @[StrongEnum.scala 204:11]
  wire  _T_983; // @[StrongEnum.scala 205:22]
  wire  _T_985; // @[StrongEnum.scala 205:11]
  wire  _T_986; // @[StrongEnum.scala 205:11]
  wire  _T_990; // @[StrongEnum.scala 206:22]
  wire  _T_992; // @[StrongEnum.scala 206:11]
  wire  _T_993; // @[StrongEnum.scala 206:11]
  wire  _T_997; // @[StrongEnum.scala 207:22]
  wire  _T_999; // @[StrongEnum.scala 207:11]
  wire  _T_1000; // @[StrongEnum.scala 207:11]
  wire  _T_1004; // @[StrongEnum.scala 208:22]
  wire  _T_1006; // @[StrongEnum.scala 208:11]
  wire  _T_1007; // @[StrongEnum.scala 208:11]
  wire  _T_1011; // @[StrongEnum.scala 203:22]
  wire  _T_1013; // @[StrongEnum.scala 203:11]
  wire  _T_1014; // @[StrongEnum.scala 203:11]
  wire  _T_1018; // @[StrongEnum.scala 204:22]
  wire  _T_1020; // @[StrongEnum.scala 204:11]
  wire  _T_1021; // @[StrongEnum.scala 204:11]
  wire  _T_1025; // @[StrongEnum.scala 205:22]
  wire  _T_1027; // @[StrongEnum.scala 205:11]
  wire  _T_1028; // @[StrongEnum.scala 205:11]
  wire  _T_1032; // @[StrongEnum.scala 206:22]
  wire  _T_1034; // @[StrongEnum.scala 206:11]
  wire  _T_1035; // @[StrongEnum.scala 206:11]
  wire  _T_1039; // @[StrongEnum.scala 207:22]
  wire  _T_1041; // @[StrongEnum.scala 207:11]
  wire  _T_1042; // @[StrongEnum.scala 207:11]
  wire  _T_1046; // @[StrongEnum.scala 208:22]
  wire  _T_1048; // @[StrongEnum.scala 208:11]
  wire  _T_1049; // @[StrongEnum.scala 208:11]
  wire  _T_1051; // @[StrongEnum.scala 210:7]
  EnumOps EnumOps ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_io_x),
    .io_y(EnumOps_io_y),
    .io_lt(EnumOps_io_lt),
    .io_le(EnumOps_io_le),
    .io_gt(EnumOps_io_gt),
    .io_ge(EnumOps_io_ge),
    .io_eq(EnumOps_io_eq),
    .io_ne(EnumOps_io_ne)
  );
  EnumOps EnumOps_1 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_1_io_x),
    .io_y(EnumOps_1_io_y),
    .io_lt(EnumOps_1_io_lt),
    .io_le(EnumOps_1_io_le),
    .io_gt(EnumOps_1_io_gt),
    .io_ge(EnumOps_1_io_ge),
    .io_eq(EnumOps_1_io_eq),
    .io_ne(EnumOps_1_io_ne)
  );
  EnumOps EnumOps_2 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_2_io_x),
    .io_y(EnumOps_2_io_y),
    .io_lt(EnumOps_2_io_lt),
    .io_le(EnumOps_2_io_le),
    .io_gt(EnumOps_2_io_gt),
    .io_ge(EnumOps_2_io_ge),
    .io_eq(EnumOps_2_io_eq),
    .io_ne(EnumOps_2_io_ne)
  );
  EnumOps EnumOps_3 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_3_io_x),
    .io_y(EnumOps_3_io_y),
    .io_lt(EnumOps_3_io_lt),
    .io_le(EnumOps_3_io_le),
    .io_gt(EnumOps_3_io_gt),
    .io_ge(EnumOps_3_io_ge),
    .io_eq(EnumOps_3_io_eq),
    .io_ne(EnumOps_3_io_ne)
  );
  EnumOps EnumOps_4 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_4_io_x),
    .io_y(EnumOps_4_io_y),
    .io_lt(EnumOps_4_io_lt),
    .io_le(EnumOps_4_io_le),
    .io_gt(EnumOps_4_io_gt),
    .io_ge(EnumOps_4_io_ge),
    .io_eq(EnumOps_4_io_eq),
    .io_ne(EnumOps_4_io_ne)
  );
  EnumOps EnumOps_5 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_5_io_x),
    .io_y(EnumOps_5_io_y),
    .io_lt(EnumOps_5_io_lt),
    .io_le(EnumOps_5_io_le),
    .io_gt(EnumOps_5_io_gt),
    .io_ge(EnumOps_5_io_ge),
    .io_eq(EnumOps_5_io_eq),
    .io_ne(EnumOps_5_io_ne)
  );
  EnumOps EnumOps_6 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_6_io_x),
    .io_y(EnumOps_6_io_y),
    .io_lt(EnumOps_6_io_lt),
    .io_le(EnumOps_6_io_le),
    .io_gt(EnumOps_6_io_gt),
    .io_ge(EnumOps_6_io_ge),
    .io_eq(EnumOps_6_io_eq),
    .io_ne(EnumOps_6_io_ne)
  );
  EnumOps EnumOps_7 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_7_io_x),
    .io_y(EnumOps_7_io_y),
    .io_lt(EnumOps_7_io_lt),
    .io_le(EnumOps_7_io_le),
    .io_gt(EnumOps_7_io_gt),
    .io_ge(EnumOps_7_io_ge),
    .io_eq(EnumOps_7_io_eq),
    .io_ne(EnumOps_7_io_ne)
  );
  EnumOps EnumOps_8 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_8_io_x),
    .io_y(EnumOps_8_io_y),
    .io_lt(EnumOps_8_io_lt),
    .io_le(EnumOps_8_io_le),
    .io_gt(EnumOps_8_io_gt),
    .io_ge(EnumOps_8_io_ge),
    .io_eq(EnumOps_8_io_eq),
    .io_ne(EnumOps_8_io_ne)
  );
  EnumOps EnumOps_9 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_9_io_x),
    .io_y(EnumOps_9_io_y),
    .io_lt(EnumOps_9_io_lt),
    .io_le(EnumOps_9_io_le),
    .io_gt(EnumOps_9_io_gt),
    .io_ge(EnumOps_9_io_ge),
    .io_eq(EnumOps_9_io_eq),
    .io_ne(EnumOps_9_io_ne)
  );
  EnumOps EnumOps_10 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_10_io_x),
    .io_y(EnumOps_10_io_y),
    .io_lt(EnumOps_10_io_lt),
    .io_le(EnumOps_10_io_le),
    .io_gt(EnumOps_10_io_gt),
    .io_ge(EnumOps_10_io_ge),
    .io_eq(EnumOps_10_io_eq),
    .io_ne(EnumOps_10_io_ne)
  );
  EnumOps EnumOps_11 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_11_io_x),
    .io_y(EnumOps_11_io_y),
    .io_lt(EnumOps_11_io_lt),
    .io_le(EnumOps_11_io_le),
    .io_gt(EnumOps_11_io_gt),
    .io_ge(EnumOps_11_io_ge),
    .io_eq(EnumOps_11_io_eq),
    .io_ne(EnumOps_11_io_ne)
  );
  EnumOps EnumOps_12 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_12_io_x),
    .io_y(EnumOps_12_io_y),
    .io_lt(EnumOps_12_io_lt),
    .io_le(EnumOps_12_io_le),
    .io_gt(EnumOps_12_io_gt),
    .io_ge(EnumOps_12_io_ge),
    .io_eq(EnumOps_12_io_eq),
    .io_ne(EnumOps_12_io_ne)
  );
  EnumOps EnumOps_13 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_13_io_x),
    .io_y(EnumOps_13_io_y),
    .io_lt(EnumOps_13_io_lt),
    .io_le(EnumOps_13_io_le),
    .io_gt(EnumOps_13_io_gt),
    .io_ge(EnumOps_13_io_ge),
    .io_eq(EnumOps_13_io_eq),
    .io_ne(EnumOps_13_io_ne)
  );
  EnumOps EnumOps_14 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_14_io_x),
    .io_y(EnumOps_14_io_y),
    .io_lt(EnumOps_14_io_lt),
    .io_le(EnumOps_14_io_le),
    .io_gt(EnumOps_14_io_gt),
    .io_ge(EnumOps_14_io_ge),
    .io_eq(EnumOps_14_io_eq),
    .io_ne(EnumOps_14_io_ne)
  );
  EnumOps EnumOps_15 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_15_io_x),
    .io_y(EnumOps_15_io_y),
    .io_lt(EnumOps_15_io_lt),
    .io_le(EnumOps_15_io_le),
    .io_gt(EnumOps_15_io_gt),
    .io_ge(EnumOps_15_io_ge),
    .io_eq(EnumOps_15_io_eq),
    .io_ne(EnumOps_15_io_ne)
  );
  EnumOps EnumOps_16 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_16_io_x),
    .io_y(EnumOps_16_io_y),
    .io_lt(EnumOps_16_io_lt),
    .io_le(EnumOps_16_io_le),
    .io_gt(EnumOps_16_io_gt),
    .io_ge(EnumOps_16_io_ge),
    .io_eq(EnumOps_16_io_eq),
    .io_ne(EnumOps_16_io_ne)
  );
  EnumOps EnumOps_17 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_17_io_x),
    .io_y(EnumOps_17_io_y),
    .io_lt(EnumOps_17_io_lt),
    .io_le(EnumOps_17_io_le),
    .io_gt(EnumOps_17_io_gt),
    .io_ge(EnumOps_17_io_ge),
    .io_eq(EnumOps_17_io_eq),
    .io_ne(EnumOps_17_io_ne)
  );
  EnumOps EnumOps_18 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_18_io_x),
    .io_y(EnumOps_18_io_y),
    .io_lt(EnumOps_18_io_lt),
    .io_le(EnumOps_18_io_le),
    .io_gt(EnumOps_18_io_gt),
    .io_ge(EnumOps_18_io_ge),
    .io_eq(EnumOps_18_io_eq),
    .io_ne(EnumOps_18_io_ne)
  );
  EnumOps EnumOps_19 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_19_io_x),
    .io_y(EnumOps_19_io_y),
    .io_lt(EnumOps_19_io_lt),
    .io_le(EnumOps_19_io_le),
    .io_gt(EnumOps_19_io_gt),
    .io_ge(EnumOps_19_io_ge),
    .io_eq(EnumOps_19_io_eq),
    .io_ne(EnumOps_19_io_ne)
  );
  EnumOps EnumOps_20 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_20_io_x),
    .io_y(EnumOps_20_io_y),
    .io_lt(EnumOps_20_io_lt),
    .io_le(EnumOps_20_io_le),
    .io_gt(EnumOps_20_io_gt),
    .io_ge(EnumOps_20_io_ge),
    .io_eq(EnumOps_20_io_eq),
    .io_ne(EnumOps_20_io_ne)
  );
  EnumOps EnumOps_21 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_21_io_x),
    .io_y(EnumOps_21_io_y),
    .io_lt(EnumOps_21_io_lt),
    .io_le(EnumOps_21_io_le),
    .io_gt(EnumOps_21_io_gt),
    .io_ge(EnumOps_21_io_ge),
    .io_eq(EnumOps_21_io_eq),
    .io_ne(EnumOps_21_io_ne)
  );
  EnumOps EnumOps_22 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_22_io_x),
    .io_y(EnumOps_22_io_y),
    .io_lt(EnumOps_22_io_lt),
    .io_le(EnumOps_22_io_le),
    .io_gt(EnumOps_22_io_gt),
    .io_ge(EnumOps_22_io_ge),
    .io_eq(EnumOps_22_io_eq),
    .io_ne(EnumOps_22_io_ne)
  );
  EnumOps EnumOps_23 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_23_io_x),
    .io_y(EnumOps_23_io_y),
    .io_lt(EnumOps_23_io_lt),
    .io_le(EnumOps_23_io_le),
    .io_gt(EnumOps_23_io_gt),
    .io_ge(EnumOps_23_io_ge),
    .io_eq(EnumOps_23_io_eq),
    .io_ne(EnumOps_23_io_ne)
  );
  EnumOps EnumOps_24 ( // @[StrongEnum.scala 199:21]
    .io_x(EnumOps_24_io_x),
    .io_y(EnumOps_24_io_y),
    .io_lt(EnumOps_24_io_lt),
    .io_le(EnumOps_24_io_le),
    .io_gt(EnumOps_24_io_gt),
    .io_ge(EnumOps_24_io_ge),
    .io_eq(EnumOps_24_io_eq),
    .io_ne(EnumOps_24_io_ne)
  );
  assign _T_3 = EnumOps_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_5 = _T_3 | reset; // @[StrongEnum.scala 203:11]
  assign _T_6 = _T_5 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_10 = EnumOps_io_le; // @[StrongEnum.scala 204:22]
  assign _T_12 = _T_10 | reset; // @[StrongEnum.scala 204:11]
  assign _T_13 = _T_12 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_17 = EnumOps_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_19 = _T_17 | reset; // @[StrongEnum.scala 205:11]
  assign _T_20 = _T_19 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_24 = EnumOps_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_26 = _T_24 | reset; // @[StrongEnum.scala 206:11]
  assign _T_27 = _T_26 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_31 = EnumOps_io_eq; // @[StrongEnum.scala 207:22]
  assign _T_33 = _T_31 | reset; // @[StrongEnum.scala 207:11]
  assign _T_34 = _T_33 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_38 = EnumOps_io_ne == 1'h0; // @[StrongEnum.scala 208:22]
  assign _T_40 = _T_38 | reset; // @[StrongEnum.scala 208:11]
  assign _T_41 = _T_40 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_45 = EnumOps_1_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_47 = _T_45 | reset; // @[StrongEnum.scala 203:11]
  assign _T_48 = _T_47 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_52 = EnumOps_1_io_le; // @[StrongEnum.scala 204:22]
  assign _T_54 = _T_52 | reset; // @[StrongEnum.scala 204:11]
  assign _T_55 = _T_54 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_59 = EnumOps_1_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_61 = _T_59 | reset; // @[StrongEnum.scala 205:11]
  assign _T_62 = _T_61 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_66 = EnumOps_1_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_68 = _T_66 | reset; // @[StrongEnum.scala 206:11]
  assign _T_69 = _T_68 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_73 = EnumOps_1_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_75 = _T_73 | reset; // @[StrongEnum.scala 207:11]
  assign _T_76 = _T_75 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_80 = EnumOps_1_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_82 = _T_80 | reset; // @[StrongEnum.scala 208:11]
  assign _T_83 = _T_82 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_87 = EnumOps_2_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_89 = _T_87 | reset; // @[StrongEnum.scala 203:11]
  assign _T_90 = _T_89 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_94 = EnumOps_2_io_le; // @[StrongEnum.scala 204:22]
  assign _T_96 = _T_94 | reset; // @[StrongEnum.scala 204:11]
  assign _T_97 = _T_96 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_101 = EnumOps_2_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_103 = _T_101 | reset; // @[StrongEnum.scala 205:11]
  assign _T_104 = _T_103 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_108 = EnumOps_2_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_110 = _T_108 | reset; // @[StrongEnum.scala 206:11]
  assign _T_111 = _T_110 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_115 = EnumOps_2_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_117 = _T_115 | reset; // @[StrongEnum.scala 207:11]
  assign _T_118 = _T_117 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_122 = EnumOps_2_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_124 = _T_122 | reset; // @[StrongEnum.scala 208:11]
  assign _T_125 = _T_124 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_129 = EnumOps_3_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_131 = _T_129 | reset; // @[StrongEnum.scala 203:11]
  assign _T_132 = _T_131 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_136 = EnumOps_3_io_le; // @[StrongEnum.scala 204:22]
  assign _T_138 = _T_136 | reset; // @[StrongEnum.scala 204:11]
  assign _T_139 = _T_138 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_143 = EnumOps_3_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_145 = _T_143 | reset; // @[StrongEnum.scala 205:11]
  assign _T_146 = _T_145 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_150 = EnumOps_3_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_152 = _T_150 | reset; // @[StrongEnum.scala 206:11]
  assign _T_153 = _T_152 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_157 = EnumOps_3_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_159 = _T_157 | reset; // @[StrongEnum.scala 207:11]
  assign _T_160 = _T_159 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_164 = EnumOps_3_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_166 = _T_164 | reset; // @[StrongEnum.scala 208:11]
  assign _T_167 = _T_166 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_171 = EnumOps_4_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_173 = _T_171 | reset; // @[StrongEnum.scala 203:11]
  assign _T_174 = _T_173 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_178 = EnumOps_4_io_le; // @[StrongEnum.scala 204:22]
  assign _T_180 = _T_178 | reset; // @[StrongEnum.scala 204:11]
  assign _T_181 = _T_180 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_185 = EnumOps_4_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_187 = _T_185 | reset; // @[StrongEnum.scala 205:11]
  assign _T_188 = _T_187 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_192 = EnumOps_4_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_194 = _T_192 | reset; // @[StrongEnum.scala 206:11]
  assign _T_195 = _T_194 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_199 = EnumOps_4_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_201 = _T_199 | reset; // @[StrongEnum.scala 207:11]
  assign _T_202 = _T_201 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_206 = EnumOps_4_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_208 = _T_206 | reset; // @[StrongEnum.scala 208:11]
  assign _T_209 = _T_208 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_213 = EnumOps_5_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_215 = _T_213 | reset; // @[StrongEnum.scala 203:11]
  assign _T_216 = _T_215 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_220 = EnumOps_5_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_222 = _T_220 | reset; // @[StrongEnum.scala 204:11]
  assign _T_223 = _T_222 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_227 = EnumOps_5_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_229 = _T_227 | reset; // @[StrongEnum.scala 205:11]
  assign _T_230 = _T_229 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_234 = EnumOps_5_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_236 = _T_234 | reset; // @[StrongEnum.scala 206:11]
  assign _T_237 = _T_236 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_241 = EnumOps_5_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_243 = _T_241 | reset; // @[StrongEnum.scala 207:11]
  assign _T_244 = _T_243 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_248 = EnumOps_5_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_250 = _T_248 | reset; // @[StrongEnum.scala 208:11]
  assign _T_251 = _T_250 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_255 = EnumOps_6_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_257 = _T_255 | reset; // @[StrongEnum.scala 203:11]
  assign _T_258 = _T_257 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_262 = EnumOps_6_io_le; // @[StrongEnum.scala 204:22]
  assign _T_264 = _T_262 | reset; // @[StrongEnum.scala 204:11]
  assign _T_265 = _T_264 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_269 = EnumOps_6_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_271 = _T_269 | reset; // @[StrongEnum.scala 205:11]
  assign _T_272 = _T_271 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_276 = EnumOps_6_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_278 = _T_276 | reset; // @[StrongEnum.scala 206:11]
  assign _T_279 = _T_278 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_283 = EnumOps_6_io_eq; // @[StrongEnum.scala 207:22]
  assign _T_285 = _T_283 | reset; // @[StrongEnum.scala 207:11]
  assign _T_286 = _T_285 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_290 = EnumOps_6_io_ne == 1'h0; // @[StrongEnum.scala 208:22]
  assign _T_292 = _T_290 | reset; // @[StrongEnum.scala 208:11]
  assign _T_293 = _T_292 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_297 = EnumOps_7_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_299 = _T_297 | reset; // @[StrongEnum.scala 203:11]
  assign _T_300 = _T_299 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_304 = EnumOps_7_io_le; // @[StrongEnum.scala 204:22]
  assign _T_306 = _T_304 | reset; // @[StrongEnum.scala 204:11]
  assign _T_307 = _T_306 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_311 = EnumOps_7_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_313 = _T_311 | reset; // @[StrongEnum.scala 205:11]
  assign _T_314 = _T_313 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_318 = EnumOps_7_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_320 = _T_318 | reset; // @[StrongEnum.scala 206:11]
  assign _T_321 = _T_320 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_325 = EnumOps_7_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_327 = _T_325 | reset; // @[StrongEnum.scala 207:11]
  assign _T_328 = _T_327 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_332 = EnumOps_7_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_334 = _T_332 | reset; // @[StrongEnum.scala 208:11]
  assign _T_335 = _T_334 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_339 = EnumOps_8_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_341 = _T_339 | reset; // @[StrongEnum.scala 203:11]
  assign _T_342 = _T_341 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_346 = EnumOps_8_io_le; // @[StrongEnum.scala 204:22]
  assign _T_348 = _T_346 | reset; // @[StrongEnum.scala 204:11]
  assign _T_349 = _T_348 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_353 = EnumOps_8_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_355 = _T_353 | reset; // @[StrongEnum.scala 205:11]
  assign _T_356 = _T_355 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_360 = EnumOps_8_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_362 = _T_360 | reset; // @[StrongEnum.scala 206:11]
  assign _T_363 = _T_362 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_367 = EnumOps_8_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_369 = _T_367 | reset; // @[StrongEnum.scala 207:11]
  assign _T_370 = _T_369 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_374 = EnumOps_8_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_376 = _T_374 | reset; // @[StrongEnum.scala 208:11]
  assign _T_377 = _T_376 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_381 = EnumOps_9_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_383 = _T_381 | reset; // @[StrongEnum.scala 203:11]
  assign _T_384 = _T_383 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_388 = EnumOps_9_io_le; // @[StrongEnum.scala 204:22]
  assign _T_390 = _T_388 | reset; // @[StrongEnum.scala 204:11]
  assign _T_391 = _T_390 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_395 = EnumOps_9_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_397 = _T_395 | reset; // @[StrongEnum.scala 205:11]
  assign _T_398 = _T_397 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_402 = EnumOps_9_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_404 = _T_402 | reset; // @[StrongEnum.scala 206:11]
  assign _T_405 = _T_404 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_409 = EnumOps_9_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_411 = _T_409 | reset; // @[StrongEnum.scala 207:11]
  assign _T_412 = _T_411 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_416 = EnumOps_9_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_418 = _T_416 | reset; // @[StrongEnum.scala 208:11]
  assign _T_419 = _T_418 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_423 = EnumOps_10_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_425 = _T_423 | reset; // @[StrongEnum.scala 203:11]
  assign _T_426 = _T_425 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_430 = EnumOps_10_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_432 = _T_430 | reset; // @[StrongEnum.scala 204:11]
  assign _T_433 = _T_432 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_437 = EnumOps_10_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_439 = _T_437 | reset; // @[StrongEnum.scala 205:11]
  assign _T_440 = _T_439 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_444 = EnumOps_10_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_446 = _T_444 | reset; // @[StrongEnum.scala 206:11]
  assign _T_447 = _T_446 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_451 = EnumOps_10_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_453 = _T_451 | reset; // @[StrongEnum.scala 207:11]
  assign _T_454 = _T_453 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_458 = EnumOps_10_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_460 = _T_458 | reset; // @[StrongEnum.scala 208:11]
  assign _T_461 = _T_460 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_465 = EnumOps_11_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_467 = _T_465 | reset; // @[StrongEnum.scala 203:11]
  assign _T_468 = _T_467 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_472 = EnumOps_11_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_474 = _T_472 | reset; // @[StrongEnum.scala 204:11]
  assign _T_475 = _T_474 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_479 = EnumOps_11_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_481 = _T_479 | reset; // @[StrongEnum.scala 205:11]
  assign _T_482 = _T_481 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_486 = EnumOps_11_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_488 = _T_486 | reset; // @[StrongEnum.scala 206:11]
  assign _T_489 = _T_488 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_493 = EnumOps_11_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_495 = _T_493 | reset; // @[StrongEnum.scala 207:11]
  assign _T_496 = _T_495 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_500 = EnumOps_11_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_502 = _T_500 | reset; // @[StrongEnum.scala 208:11]
  assign _T_503 = _T_502 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_507 = EnumOps_12_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_509 = _T_507 | reset; // @[StrongEnum.scala 203:11]
  assign _T_510 = _T_509 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_514 = EnumOps_12_io_le; // @[StrongEnum.scala 204:22]
  assign _T_516 = _T_514 | reset; // @[StrongEnum.scala 204:11]
  assign _T_517 = _T_516 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_521 = EnumOps_12_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_523 = _T_521 | reset; // @[StrongEnum.scala 205:11]
  assign _T_524 = _T_523 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_528 = EnumOps_12_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_530 = _T_528 | reset; // @[StrongEnum.scala 206:11]
  assign _T_531 = _T_530 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_535 = EnumOps_12_io_eq; // @[StrongEnum.scala 207:22]
  assign _T_537 = _T_535 | reset; // @[StrongEnum.scala 207:11]
  assign _T_538 = _T_537 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_542 = EnumOps_12_io_ne == 1'h0; // @[StrongEnum.scala 208:22]
  assign _T_544 = _T_542 | reset; // @[StrongEnum.scala 208:11]
  assign _T_545 = _T_544 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_549 = EnumOps_13_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_551 = _T_549 | reset; // @[StrongEnum.scala 203:11]
  assign _T_552 = _T_551 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_556 = EnumOps_13_io_le; // @[StrongEnum.scala 204:22]
  assign _T_558 = _T_556 | reset; // @[StrongEnum.scala 204:11]
  assign _T_559 = _T_558 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_563 = EnumOps_13_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_565 = _T_563 | reset; // @[StrongEnum.scala 205:11]
  assign _T_566 = _T_565 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_570 = EnumOps_13_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_572 = _T_570 | reset; // @[StrongEnum.scala 206:11]
  assign _T_573 = _T_572 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_577 = EnumOps_13_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_579 = _T_577 | reset; // @[StrongEnum.scala 207:11]
  assign _T_580 = _T_579 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_584 = EnumOps_13_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_586 = _T_584 | reset; // @[StrongEnum.scala 208:11]
  assign _T_587 = _T_586 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_591 = EnumOps_14_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_593 = _T_591 | reset; // @[StrongEnum.scala 203:11]
  assign _T_594 = _T_593 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_598 = EnumOps_14_io_le; // @[StrongEnum.scala 204:22]
  assign _T_600 = _T_598 | reset; // @[StrongEnum.scala 204:11]
  assign _T_601 = _T_600 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_605 = EnumOps_14_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_607 = _T_605 | reset; // @[StrongEnum.scala 205:11]
  assign _T_608 = _T_607 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_612 = EnumOps_14_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_614 = _T_612 | reset; // @[StrongEnum.scala 206:11]
  assign _T_615 = _T_614 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_619 = EnumOps_14_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_621 = _T_619 | reset; // @[StrongEnum.scala 207:11]
  assign _T_622 = _T_621 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_626 = EnumOps_14_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_628 = _T_626 | reset; // @[StrongEnum.scala 208:11]
  assign _T_629 = _T_628 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_633 = EnumOps_15_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_635 = _T_633 | reset; // @[StrongEnum.scala 203:11]
  assign _T_636 = _T_635 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_640 = EnumOps_15_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_642 = _T_640 | reset; // @[StrongEnum.scala 204:11]
  assign _T_643 = _T_642 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_647 = EnumOps_15_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_649 = _T_647 | reset; // @[StrongEnum.scala 205:11]
  assign _T_650 = _T_649 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_654 = EnumOps_15_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_656 = _T_654 | reset; // @[StrongEnum.scala 206:11]
  assign _T_657 = _T_656 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_661 = EnumOps_15_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_663 = _T_661 | reset; // @[StrongEnum.scala 207:11]
  assign _T_664 = _T_663 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_668 = EnumOps_15_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_670 = _T_668 | reset; // @[StrongEnum.scala 208:11]
  assign _T_671 = _T_670 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_675 = EnumOps_16_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_677 = _T_675 | reset; // @[StrongEnum.scala 203:11]
  assign _T_678 = _T_677 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_682 = EnumOps_16_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_684 = _T_682 | reset; // @[StrongEnum.scala 204:11]
  assign _T_685 = _T_684 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_689 = EnumOps_16_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_691 = _T_689 | reset; // @[StrongEnum.scala 205:11]
  assign _T_692 = _T_691 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_696 = EnumOps_16_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_698 = _T_696 | reset; // @[StrongEnum.scala 206:11]
  assign _T_699 = _T_698 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_703 = EnumOps_16_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_705 = _T_703 | reset; // @[StrongEnum.scala 207:11]
  assign _T_706 = _T_705 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_710 = EnumOps_16_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_712 = _T_710 | reset; // @[StrongEnum.scala 208:11]
  assign _T_713 = _T_712 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_717 = EnumOps_17_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_719 = _T_717 | reset; // @[StrongEnum.scala 203:11]
  assign _T_720 = _T_719 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_724 = EnumOps_17_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_726 = _T_724 | reset; // @[StrongEnum.scala 204:11]
  assign _T_727 = _T_726 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_731 = EnumOps_17_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_733 = _T_731 | reset; // @[StrongEnum.scala 205:11]
  assign _T_734 = _T_733 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_738 = EnumOps_17_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_740 = _T_738 | reset; // @[StrongEnum.scala 206:11]
  assign _T_741 = _T_740 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_745 = EnumOps_17_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_747 = _T_745 | reset; // @[StrongEnum.scala 207:11]
  assign _T_748 = _T_747 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_752 = EnumOps_17_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_754 = _T_752 | reset; // @[StrongEnum.scala 208:11]
  assign _T_755 = _T_754 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_759 = EnumOps_18_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_761 = _T_759 | reset; // @[StrongEnum.scala 203:11]
  assign _T_762 = _T_761 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_766 = EnumOps_18_io_le; // @[StrongEnum.scala 204:22]
  assign _T_768 = _T_766 | reset; // @[StrongEnum.scala 204:11]
  assign _T_769 = _T_768 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_773 = EnumOps_18_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_775 = _T_773 | reset; // @[StrongEnum.scala 205:11]
  assign _T_776 = _T_775 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_780 = EnumOps_18_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_782 = _T_780 | reset; // @[StrongEnum.scala 206:11]
  assign _T_783 = _T_782 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_787 = EnumOps_18_io_eq; // @[StrongEnum.scala 207:22]
  assign _T_789 = _T_787 | reset; // @[StrongEnum.scala 207:11]
  assign _T_790 = _T_789 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_794 = EnumOps_18_io_ne == 1'h0; // @[StrongEnum.scala 208:22]
  assign _T_796 = _T_794 | reset; // @[StrongEnum.scala 208:11]
  assign _T_797 = _T_796 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_801 = EnumOps_19_io_lt; // @[StrongEnum.scala 203:22]
  assign _T_803 = _T_801 | reset; // @[StrongEnum.scala 203:11]
  assign _T_804 = _T_803 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_808 = EnumOps_19_io_le; // @[StrongEnum.scala 204:22]
  assign _T_810 = _T_808 | reset; // @[StrongEnum.scala 204:11]
  assign _T_811 = _T_810 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_815 = EnumOps_19_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_817 = _T_815 | reset; // @[StrongEnum.scala 205:11]
  assign _T_818 = _T_817 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_822 = EnumOps_19_io_ge == 1'h0; // @[StrongEnum.scala 206:22]
  assign _T_824 = _T_822 | reset; // @[StrongEnum.scala 206:11]
  assign _T_825 = _T_824 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_829 = EnumOps_19_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_831 = _T_829 | reset; // @[StrongEnum.scala 207:11]
  assign _T_832 = _T_831 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_836 = EnumOps_19_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_838 = _T_836 | reset; // @[StrongEnum.scala 208:11]
  assign _T_839 = _T_838 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_843 = EnumOps_20_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_845 = _T_843 | reset; // @[StrongEnum.scala 203:11]
  assign _T_846 = _T_845 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_850 = EnumOps_20_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_852 = _T_850 | reset; // @[StrongEnum.scala 204:11]
  assign _T_853 = _T_852 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_857 = EnumOps_20_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_859 = _T_857 | reset; // @[StrongEnum.scala 205:11]
  assign _T_860 = _T_859 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_864 = EnumOps_20_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_866 = _T_864 | reset; // @[StrongEnum.scala 206:11]
  assign _T_867 = _T_866 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_871 = EnumOps_20_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_873 = _T_871 | reset; // @[StrongEnum.scala 207:11]
  assign _T_874 = _T_873 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_878 = EnumOps_20_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_880 = _T_878 | reset; // @[StrongEnum.scala 208:11]
  assign _T_881 = _T_880 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_885 = EnumOps_21_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_887 = _T_885 | reset; // @[StrongEnum.scala 203:11]
  assign _T_888 = _T_887 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_892 = EnumOps_21_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_894 = _T_892 | reset; // @[StrongEnum.scala 204:11]
  assign _T_895 = _T_894 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_899 = EnumOps_21_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_901 = _T_899 | reset; // @[StrongEnum.scala 205:11]
  assign _T_902 = _T_901 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_906 = EnumOps_21_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_908 = _T_906 | reset; // @[StrongEnum.scala 206:11]
  assign _T_909 = _T_908 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_913 = EnumOps_21_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_915 = _T_913 | reset; // @[StrongEnum.scala 207:11]
  assign _T_916 = _T_915 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_920 = EnumOps_21_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_922 = _T_920 | reset; // @[StrongEnum.scala 208:11]
  assign _T_923 = _T_922 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_927 = EnumOps_22_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_929 = _T_927 | reset; // @[StrongEnum.scala 203:11]
  assign _T_930 = _T_929 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_934 = EnumOps_22_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_936 = _T_934 | reset; // @[StrongEnum.scala 204:11]
  assign _T_937 = _T_936 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_941 = EnumOps_22_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_943 = _T_941 | reset; // @[StrongEnum.scala 205:11]
  assign _T_944 = _T_943 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_948 = EnumOps_22_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_950 = _T_948 | reset; // @[StrongEnum.scala 206:11]
  assign _T_951 = _T_950 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_955 = EnumOps_22_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_957 = _T_955 | reset; // @[StrongEnum.scala 207:11]
  assign _T_958 = _T_957 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_962 = EnumOps_22_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_964 = _T_962 | reset; // @[StrongEnum.scala 208:11]
  assign _T_965 = _T_964 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_969 = EnumOps_23_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_971 = _T_969 | reset; // @[StrongEnum.scala 203:11]
  assign _T_972 = _T_971 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_976 = EnumOps_23_io_le == 1'h0; // @[StrongEnum.scala 204:22]
  assign _T_978 = _T_976 | reset; // @[StrongEnum.scala 204:11]
  assign _T_979 = _T_978 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_983 = EnumOps_23_io_gt; // @[StrongEnum.scala 205:22]
  assign _T_985 = _T_983 | reset; // @[StrongEnum.scala 205:11]
  assign _T_986 = _T_985 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_990 = EnumOps_23_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_992 = _T_990 | reset; // @[StrongEnum.scala 206:11]
  assign _T_993 = _T_992 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_997 = EnumOps_23_io_eq == 1'h0; // @[StrongEnum.scala 207:22]
  assign _T_999 = _T_997 | reset; // @[StrongEnum.scala 207:11]
  assign _T_1000 = _T_999 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_1004 = EnumOps_23_io_ne; // @[StrongEnum.scala 208:22]
  assign _T_1006 = _T_1004 | reset; // @[StrongEnum.scala 208:11]
  assign _T_1007 = _T_1006 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_1011 = EnumOps_24_io_lt == 1'h0; // @[StrongEnum.scala 203:22]
  assign _T_1013 = _T_1011 | reset; // @[StrongEnum.scala 203:11]
  assign _T_1014 = _T_1013 == 1'h0; // @[StrongEnum.scala 203:11]
  assign _T_1018 = EnumOps_24_io_le; // @[StrongEnum.scala 204:22]
  assign _T_1020 = _T_1018 | reset; // @[StrongEnum.scala 204:11]
  assign _T_1021 = _T_1020 == 1'h0; // @[StrongEnum.scala 204:11]
  assign _T_1025 = EnumOps_24_io_gt == 1'h0; // @[StrongEnum.scala 205:22]
  assign _T_1027 = _T_1025 | reset; // @[StrongEnum.scala 205:11]
  assign _T_1028 = _T_1027 == 1'h0; // @[StrongEnum.scala 205:11]
  assign _T_1032 = EnumOps_24_io_ge; // @[StrongEnum.scala 206:22]
  assign _T_1034 = _T_1032 | reset; // @[StrongEnum.scala 206:11]
  assign _T_1035 = _T_1034 == 1'h0; // @[StrongEnum.scala 206:11]
  assign _T_1039 = EnumOps_24_io_eq; // @[StrongEnum.scala 207:22]
  assign _T_1041 = _T_1039 | reset; // @[StrongEnum.scala 207:11]
  assign _T_1042 = _T_1041 == 1'h0; // @[StrongEnum.scala 207:11]
  assign _T_1046 = EnumOps_24_io_ne == 1'h0; // @[StrongEnum.scala 208:22]
  assign _T_1048 = _T_1046 | reset; // @[StrongEnum.scala 208:11]
  assign _T_1049 = _T_1048 == 1'h0; // @[StrongEnum.scala 208:11]
  assign _T_1051 = reset == 1'h0; // @[StrongEnum.scala 210:7]
  assign EnumOps_io_x = 7'h0; // @[StrongEnum.scala 200:14]
  assign EnumOps_io_y = 7'h0; // @[StrongEnum.scala 201:14]
  assign EnumOps_1_io_x = 7'h0; // @[StrongEnum.scala 200:14]
  assign EnumOps_1_io_y = 7'h1; // @[StrongEnum.scala 201:14]
  assign EnumOps_2_io_x = 7'h0; // @[StrongEnum.scala 200:14]
  assign EnumOps_2_io_y = 7'h2; // @[StrongEnum.scala 201:14]
  assign EnumOps_3_io_x = 7'h0; // @[StrongEnum.scala 200:14]
  assign EnumOps_3_io_y = 7'h64; // @[StrongEnum.scala 201:14]
  assign EnumOps_4_io_x = 7'h0; // @[StrongEnum.scala 200:14]
  assign EnumOps_4_io_y = 7'h65; // @[StrongEnum.scala 201:14]
  assign EnumOps_5_io_x = 7'h1; // @[StrongEnum.scala 200:14]
  assign EnumOps_5_io_y = 7'h0; // @[StrongEnum.scala 201:14]
  assign EnumOps_6_io_x = 7'h1; // @[StrongEnum.scala 200:14]
  assign EnumOps_6_io_y = 7'h1; // @[StrongEnum.scala 201:14]
  assign EnumOps_7_io_x = 7'h1; // @[StrongEnum.scala 200:14]
  assign EnumOps_7_io_y = 7'h2; // @[StrongEnum.scala 201:14]
  assign EnumOps_8_io_x = 7'h1; // @[StrongEnum.scala 200:14]
  assign EnumOps_8_io_y = 7'h64; // @[StrongEnum.scala 201:14]
  assign EnumOps_9_io_x = 7'h1; // @[StrongEnum.scala 200:14]
  assign EnumOps_9_io_y = 7'h65; // @[StrongEnum.scala 201:14]
  assign EnumOps_10_io_x = 7'h2; // @[StrongEnum.scala 200:14]
  assign EnumOps_10_io_y = 7'h0; // @[StrongEnum.scala 201:14]
  assign EnumOps_11_io_x = 7'h2; // @[StrongEnum.scala 200:14]
  assign EnumOps_11_io_y = 7'h1; // @[StrongEnum.scala 201:14]
  assign EnumOps_12_io_x = 7'h2; // @[StrongEnum.scala 200:14]
  assign EnumOps_12_io_y = 7'h2; // @[StrongEnum.scala 201:14]
  assign EnumOps_13_io_x = 7'h2; // @[StrongEnum.scala 200:14]
  assign EnumOps_13_io_y = 7'h64; // @[StrongEnum.scala 201:14]
  assign EnumOps_14_io_x = 7'h2; // @[StrongEnum.scala 200:14]
  assign EnumOps_14_io_y = 7'h65; // @[StrongEnum.scala 201:14]
  assign EnumOps_15_io_x = 7'h64; // @[StrongEnum.scala 200:14]
  assign EnumOps_15_io_y = 7'h0; // @[StrongEnum.scala 201:14]
  assign EnumOps_16_io_x = 7'h64; // @[StrongEnum.scala 200:14]
  assign EnumOps_16_io_y = 7'h1; // @[StrongEnum.scala 201:14]
  assign EnumOps_17_io_x = 7'h64; // @[StrongEnum.scala 200:14]
  assign EnumOps_17_io_y = 7'h2; // @[StrongEnum.scala 201:14]
  assign EnumOps_18_io_x = 7'h64; // @[StrongEnum.scala 200:14]
  assign EnumOps_18_io_y = 7'h64; // @[StrongEnum.scala 201:14]
  assign EnumOps_19_io_x = 7'h64; // @[StrongEnum.scala 200:14]
  assign EnumOps_19_io_y = 7'h65; // @[StrongEnum.scala 201:14]
  assign EnumOps_20_io_x = 7'h65; // @[StrongEnum.scala 200:14]
  assign EnumOps_20_io_y = 7'h0; // @[StrongEnum.scala 201:14]
  assign EnumOps_21_io_x = 7'h65; // @[StrongEnum.scala 200:14]
  assign EnumOps_21_io_y = 7'h1; // @[StrongEnum.scala 201:14]
  assign EnumOps_22_io_x = 7'h65; // @[StrongEnum.scala 200:14]
  assign EnumOps_22_io_y = 7'h2; // @[StrongEnum.scala 201:14]
  assign EnumOps_23_io_x = 7'h65; // @[StrongEnum.scala 200:14]
  assign EnumOps_23_io_y = 7'h64; // @[StrongEnum.scala 201:14]
  assign EnumOps_24_io_x = 7'h65; // @[StrongEnum.scala 200:14]
  assign EnumOps_24_io_y = 7'h65; // @[StrongEnum.scala 201:14]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_20) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_27) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_27) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_34) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_34) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_41) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_48) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_48) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_55) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_55) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_62) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_62) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_69) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_69) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_76) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_76) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_83) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_83) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_90) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_90) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_97) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_97) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_104) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_111) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_111) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_118) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_118) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_125) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_125) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_132) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_132) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_139) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_139) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_146) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_146) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_153) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_153) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_160) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_160) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_167) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_167) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_174) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_174) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_181) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_181) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_188) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_188) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_195) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_195) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_202) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_202) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_209) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_209) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_216) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_216) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_223) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_223) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_230) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_230) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_237) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_237) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_244) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_244) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_251) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_251) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_258) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_258) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_265) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_265) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_272) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_272) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_279) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_279) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_286) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_286) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_293) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_293) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_300) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_300) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_307) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_307) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_314) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_314) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_321) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_321) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_328) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_328) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_335) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_335) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_342) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_342) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_349) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_349) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_356) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_356) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_363) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_363) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_370) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_370) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_377) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_377) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_384) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_384) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_391) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_391) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_398) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_398) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_405) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_405) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_412) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_412) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_419) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_419) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_426) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_426) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_433) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_433) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_440) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_440) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_447) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_447) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_454) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_454) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_461) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_461) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_468) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_468) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_475) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_475) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_482) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_482) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_489) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_489) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_496) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_496) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_503) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_503) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_510) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_510) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_517) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_517) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_524) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_524) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_531) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_531) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_538) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_538) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_545) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_545) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_559) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_559) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_566) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_566) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_573) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_573) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_580) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_580) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_587) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_587) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_594) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_594) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_615) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_615) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_622) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_622) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_629) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_629) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_636) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_636) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_643) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_643) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_650) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_650) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_657) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_657) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_671) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_671) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_678) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_678) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_685) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_685) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_692) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_692) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_706) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_706) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_713) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_713) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_720) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_720) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_727) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_727) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_734) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_734) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_741) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_741) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_748) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_748) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_755) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_755) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_762) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_762) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_769) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_769) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_776) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_776) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_783) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_783) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_790) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_790) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_797) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_797) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_804) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_804) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_811) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_811) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_818) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_818) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_825) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_825) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_839) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_839) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_846) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_846) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_853) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_853) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_860) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_860) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_867) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_867) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_874) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_874) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_881) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_881) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_888) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_888) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_895) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_895) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_902) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_902) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_909) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_909) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_916) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_916) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_923) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_923) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_930) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_930) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_937) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_937) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_944) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_944) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_951) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_951) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_958) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_958) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_965) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_965) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_972) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_972) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_979) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_979) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_986) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_986) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_993) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_993) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1000) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1000) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1007) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1007) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1014) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:203 assert(mod.io.lt === (x.asUInt() < y.asUInt()))\n"); // @[StrongEnum.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1014) begin
          $fatal; // @[StrongEnum.scala 203:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1021) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:204 assert(mod.io.le === (x.asUInt() <= y.asUInt()))\n"); // @[StrongEnum.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1021) begin
          $fatal; // @[StrongEnum.scala 204:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1028) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:205 assert(mod.io.gt === (x.asUInt() > y.asUInt()))\n"); // @[StrongEnum.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1028) begin
          $fatal; // @[StrongEnum.scala 205:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1035) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:206 assert(mod.io.ge === (x.asUInt() >= y.asUInt()))\n"); // @[StrongEnum.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1035) begin
          $fatal; // @[StrongEnum.scala 206:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1042) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:207 assert(mod.io.eq === (x.asUInt() === y.asUInt()))\n"); // @[StrongEnum.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1042) begin
          $fatal; // @[StrongEnum.scala 207:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1049) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:208 assert(mod.io.ne === (x.asUInt() =/= y.asUInt()))\n"); // @[StrongEnum.scala 208:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1049) begin
          $fatal; // @[StrongEnum.scala 208:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1051) begin
          $finish; // @[StrongEnum.scala 210:7]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
