module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [6:0]  io_in_sExp,
  input  [11:0] io_in_sig,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire [8:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [9:0] _T_3; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [9:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire [26:0] adjustedSig; // @[RoundAnyRawFNToRecFN.scala 112:22]
  wire [9:0] _T_6; // @[RoundAnyRawFNToRecFN.scala 134:55]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 134:55]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 138:28]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire [8:0] _T_22; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_24; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_32; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_34; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_39; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_41; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_42; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire [22:0] _T_44; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] _T_48; // @[Cat.scala 29:58]
  wire [2:0] _T_52; // @[Cat.scala 29:58]
  assign _GEN_0 = {{2{io_in_sExp[6]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign _T_3 = $signed(_GEN_0) + 9'she0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_T_3[8:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign adjustedSig = {io_in_sig, 15'h0}; // @[RoundAnyRawFNToRecFN.scala 112:22]
  assign _T_6 = {{1'd0}, sAdjustedExp[8:0]}; // @[RoundAnyRawFNToRecFN.scala 134:55]
  assign common_expOut = _T_6[8:0]; // @[RoundAnyRawFNToRecFN.scala 134:55]
  assign common_fractOut = adjustedSig[24:2]; // @[RoundAnyRawFNToRecFN.scala 138:28]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_22 = io_in_isZero ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_24 = common_expOut & ~_T_22; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_32 = io_in_isInf ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_34 = _T_24 & ~_T_32; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_39 = io_in_isInf ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_40 = _T_34 | _T_39; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_41 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_40 | _T_41; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_42 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_44 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign fractOut = _T_42 ? _T_44 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_48 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_52 = {io_invalidExc,1'h0,1'h0}; // @[Cat.scala 29:58]
  assign io_out = {_T_48,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_52,2'h0}; // @[RoundAnyRawFNToRecFN.scala 285:23]
endmodule
module RecFNToRecFN(
  input  [16:0] io_in,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  RoundAnyRawFNToRecFN_io_invalidExc; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isNaN; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isInf; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isZero; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_sign; // @[RecFNToRecFN.scala 72:19]
  wire [6:0] RoundAnyRawFNToRecFN_io_in_sExp; // @[RecFNToRecFN.scala 72:19]
  wire [11:0] RoundAnyRawFNToRecFN_io_in_sig; // @[RecFNToRecFN.scala 72:19]
  wire [32:0] RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 72:19]
  wire [4:0] RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 72:19]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [11:0] rawIn_sig; // @[Cat.scala 29:58]
  RoundAnyRawFNToRecFN RoundAnyRawFNToRecFN ( // @[RecFNToRecFN.scala 72:19]
    .io_invalidExc(RoundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(RoundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(RoundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(RoundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(RoundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(RoundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(RoundAnyRawFNToRecFN_io_in_sig),
    .io_out(RoundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(RoundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign rawIn_isZero = io_in[15:13] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_in[15:14] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_4 & io_in[13]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_14 = {1'h0,~rawIn_isZero}; // @[Cat.scala 29:58]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[9:0]}; // @[Cat.scala 29:58]
  assign io_out = RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 85:27]
  assign io_exceptionFlags = RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 86:27]
  assign RoundAnyRawFNToRecFN_io_invalidExc = rawIn_isNaN & ~rawIn_sig[9]; // @[RecFNToRecFN.scala 80:48]
  assign RoundAnyRawFNToRecFN_io_in_isNaN = _T_4 & io_in[13]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isInf = _T_4 & ~io_in[13]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isZero = io_in[15:13] == 3'h0; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sign = io_in[16]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(io_in[15:10])}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sig = {_T_14,io_in[9:0]}; // @[RecFNToRecFN.scala 82:48]
endmodule
module ValExec_RecF16ToRecF32(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [31:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [32:0] io_expected_recOut,
  output [32:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [16:0] recFNToRecFN_io_in; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire [32:0] recFNToRecFN_io_out; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire [4:0] recFNToRecFN_io_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_15; // @[Mux.scala 47:69]
  wire [3:0] _T_16; // @[Mux.scala 47:69]
  wire [3:0] _T_17; // @[Mux.scala 47:69]
  wire [3:0] _T_18; // @[Mux.scala 47:69]
  wire [3:0] _T_19; // @[Mux.scala 47:69]
  wire [3:0] _T_20; // @[Mux.scala 47:69]
  wire [3:0] _T_21; // @[Mux.scala 47:69]
  wire [3:0] _T_22; // @[Mux.scala 47:69]
  wire [3:0] _T_23; // @[Mux.scala 47:69]
  wire [24:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_24; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_26; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_27; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_28; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_29; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_30; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_32; // @[rawFloatFromFN.scala 59:15]
  wire  _T_33; // @[rawFloatFromFN.scala 62:34]
  wire  _T_35; // @[rawFloatFromFN.scala 63:62]
  wire  _T_38; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_41; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_43; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_45; // @[Cat.scala 29:58]
  wire [2:0] _T_47; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_49; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_52; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[Cat.scala 29:58]
  wire  _T_58; // @[rawFloatFromFN.scala 50:34]
  wire  _T_59; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_83; // @[Mux.scala 47:69]
  wire [4:0] _T_84; // @[Mux.scala 47:69]
  wire [4:0] _T_85; // @[Mux.scala 47:69]
  wire [4:0] _T_86; // @[Mux.scala 47:69]
  wire [4:0] _T_87; // @[Mux.scala 47:69]
  wire [4:0] _T_88; // @[Mux.scala 47:69]
  wire [4:0] _T_89; // @[Mux.scala 47:69]
  wire [4:0] _T_90; // @[Mux.scala 47:69]
  wire [4:0] _T_91; // @[Mux.scala 47:69]
  wire [4:0] _T_92; // @[Mux.scala 47:69]
  wire [4:0] _T_93; // @[Mux.scala 47:69]
  wire [4:0] _T_94; // @[Mux.scala 47:69]
  wire [4:0] _T_95; // @[Mux.scala 47:69]
  wire [4:0] _T_96; // @[Mux.scala 47:69]
  wire [4:0] _T_97; // @[Mux.scala 47:69]
  wire [4:0] _T_98; // @[Mux.scala 47:69]
  wire [4:0] _T_99; // @[Mux.scala 47:69]
  wire [4:0] _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_104; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_105; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_107; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_108; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_109; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_110; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_111; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_113; // @[rawFloatFromFN.scala 59:15]
  wire  _T_114; // @[rawFloatFromFN.scala 62:34]
  wire  _T_116; // @[rawFloatFromFN.scala 63:62]
  wire  _T_119; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_122; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_124; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_126; // @[Cat.scala 29:58]
  wire [2:0] _T_128; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_130; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_133; // @[Cat.scala 29:58]
  wire [3:0] _T_134; // @[Cat.scala 29:58]
  wire  _T_139; // @[tests.scala 48:26]
  wire  _T_141; // @[tests.scala 48:55]
  wire  _T_142; // @[tests.scala 48:39]
  wire  _T_143; // @[tests.scala 49:20]
  wire  _T_146; // @[tests.scala 49:54]
  wire  _T_147; // @[tests.scala 49:31]
  wire  _T_149; // @[tests.scala 50:30]
  wire  _T_151; // @[tests.scala 50:66]
  wire  _T_152; // @[tests.scala 50:16]
  wire  _T_153; // @[tests.scala 48:12]
  wire  _T_154; // @[ValExec_RecFNToRecFN.scala 84:35]
  RecFNToRecFN recFNToRecFN ( // @[ValExec_RecFNToRecFN.scala 68:15]
    .io_in(recFNToRecFN_io_in),
    .io_out(recFNToRecFN_io_out),
    .io_exceptionFlags(recFNToRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_in[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_in[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_15 = io_in[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_16 = io_in[2] ? 4'h7 : _T_15; // @[Mux.scala 47:69]
  assign _T_17 = io_in[3] ? 4'h6 : _T_16; // @[Mux.scala 47:69]
  assign _T_18 = io_in[4] ? 4'h5 : _T_17; // @[Mux.scala 47:69]
  assign _T_19 = io_in[5] ? 4'h4 : _T_18; // @[Mux.scala 47:69]
  assign _T_20 = io_in[6] ? 4'h3 : _T_19; // @[Mux.scala 47:69]
  assign _T_21 = io_in[7] ? 4'h2 : _T_20; // @[Mux.scala 47:69]
  assign _T_22 = io_in[8] ? 4'h1 : _T_21; // @[Mux.scala 47:69]
  assign _T_23 = io_in[9] ? 4'h0 : _T_22; // @[Mux.scala 47:69]
  assign _GEN_0 = {{15'd0}, io_in[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_24 = _GEN_0 << _T_23; // @[rawFloatFromFN.scala 54:36]
  assign _T_26 = {_T_24[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{2'd0}, _T_23}; // @[rawFloatFromFN.scala 57:26]
  assign _T_27 = _GEN_1 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_28 = _T_3 ? _T_27 : {{1'd0}, io_in[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_29 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{3'd0}, _T_29}; // @[rawFloatFromFN.scala 60:22]
  assign _T_30 = 5'h10 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_30}; // @[rawFloatFromFN.scala 59:15]
  assign _T_32 = _T_28 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_33 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_35 = _T_32[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_38 = _T_35 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_41 = {1'b0,$signed(_T_32)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_43 = _T_3 ? _T_26 : io_in[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_45 = {1'h0,~_T_33,_T_43}; // @[Cat.scala 29:58]
  assign _T_47 = _T_33 ? 3'h0 : _T_41[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_38}; // @[recFNFromFN.scala 48:79]
  assign _T_49 = _T_47 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_52 = {_T_41[2:0],_T_45[9:0]}; // @[Cat.scala 29:58]
  assign _T_53 = {io_in[15],_T_49}; // @[Cat.scala 29:58]
  assign _T_58 = io_expected_out[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_59 = io_expected_out[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_83 = io_expected_out[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_84 = io_expected_out[2] ? 5'h14 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = io_expected_out[3] ? 5'h13 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = io_expected_out[4] ? 5'h12 : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = io_expected_out[5] ? 5'h11 : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = io_expected_out[6] ? 5'h10 : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = io_expected_out[7] ? 5'hf : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = io_expected_out[8] ? 5'he : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = io_expected_out[9] ? 5'hd : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = io_expected_out[10] ? 5'hc : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = io_expected_out[11] ? 5'hb : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = io_expected_out[12] ? 5'ha : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = io_expected_out[13] ? 5'h9 : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = io_expected_out[14] ? 5'h8 : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = io_expected_out[15] ? 5'h7 : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = io_expected_out[16] ? 5'h6 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = io_expected_out[17] ? 5'h5 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = io_expected_out[18] ? 5'h4 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = io_expected_out[19] ? 5'h3 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = io_expected_out[20] ? 5'h2 : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = io_expected_out[21] ? 5'h1 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = io_expected_out[22] ? 5'h0 : _T_103; // @[Mux.scala 47:69]
  assign _GEN_5 = {{31'd0}, io_expected_out[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_105 = _GEN_5 << _T_104; // @[rawFloatFromFN.scala 54:36]
  assign _T_107 = {_T_105[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{4'd0}, _T_104}; // @[rawFloatFromFN.scala 57:26]
  assign _T_108 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_109 = _T_58 ? _T_108 : {{1'd0}, io_expected_out[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_110 = _T_58 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{6'd0}, _T_110}; // @[rawFloatFromFN.scala 60:22]
  assign _T_111 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_111}; // @[rawFloatFromFN.scala 59:15]
  assign _T_113 = _T_109 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_114 = _T_58 & _T_59; // @[rawFloatFromFN.scala 62:34]
  assign _T_116 = _T_113[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_119 = _T_116 & ~_T_59; // @[rawFloatFromFN.scala 66:33]
  assign _T_122 = {1'b0,$signed(_T_113)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_124 = _T_58 ? _T_107 : io_expected_out[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_126 = {1'h0,~_T_114,_T_124}; // @[Cat.scala 29:58]
  assign _T_128 = _T_114 ? 3'h0 : _T_122[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_119}; // @[recFNFromFN.scala 48:79]
  assign _T_130 = _T_128 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_133 = {_T_122[5:0],_T_126[22:0]}; // @[Cat.scala 29:58]
  assign _T_134 = {io_expected_out[31],_T_130}; // @[Cat.scala 29:58]
  assign _T_139 = io_actual_out[31:29] == 3'h0; // @[tests.scala 48:26]
  assign _T_141 = io_actual_out[31:29] == 3'h7; // @[tests.scala 48:55]
  assign _T_142 = _T_139 | _T_141; // @[tests.scala 48:39]
  assign _T_143 = io_actual_out[32:29] == io_expected_recOut[32:29]; // @[tests.scala 49:20]
  assign _T_146 = io_actual_out[22:0] == io_expected_recOut[22:0]; // @[tests.scala 49:54]
  assign _T_147 = _T_143 & _T_146; // @[tests.scala 49:31]
  assign _T_149 = io_actual_out[31:29] == 3'h6; // @[tests.scala 50:30]
  assign _T_151 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_152 = _T_149 ? _T_143 : _T_151; // @[tests.scala 50:16]
  assign _T_153 = _T_142 ? _T_147 : _T_152; // @[tests.scala 48:12]
  assign _T_154 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 84:35]
  assign io_expected_recOut = {_T_134,_T_133}; // @[ValExec_RecFNToRecFN.scala 74:24]
  assign io_actual_out = recFNToRecFN_io_out; // @[ValExec_RecFNToRecFN.scala 77:19]
  assign io_actual_exceptionFlags = recFNToRecFN_io_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 78:30]
  assign io_check = 1'h1; // @[ValExec_RecFNToRecFN.scala 80:14]
  assign io_pass = _T_153 & _T_154; // @[ValExec_RecFNToRecFN.scala 81:13]
  assign recFNToRecFN_io_in = {_T_53,_T_52}; // @[ValExec_RecFNToRecFN.scala 70:24]
endmodule
