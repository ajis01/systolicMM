module MulAddRecFNToRaw_preMul(
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [9:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [4:0]  io_toPostMul_CDom_CAlignDist,
  output [25:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawB_sig; // @[Cat.scala 29:58]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_36; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawC_sig; // @[Cat.scala 29:58]
  wire  signProd; // @[MulAddRecFN.scala 98:30]
  wire [10:0] _T_50; // @[MulAddRecFN.scala 101:19]
  wire [10:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  doSubMags; // @[MulAddRecFN.scala 103:30]
  wire [10:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [10:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [9:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _T_57; // @[MulAddRecFN.scala 109:35]
  wire  _T_58; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _T_60; // @[MulAddRecFN.scala 111:60]
  wire  _T_61; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _T_62; // @[MulAddRecFN.scala 115:34]
  wire [6:0] _T_64; // @[MulAddRecFN.scala 115:16]
  wire [6:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [24:0] _T_66; // @[MulAddRecFN.scala 121:16]
  wire [52:0] _T_68; // @[Bitwise.scala 71:12]
  wire [77:0] _T_70; // @[MulAddRecFN.scala 123:11]
  wire [77:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire [26:0] _T_71; // @[MulAddRecFN.scala 125:30]
  wire  _T_74; // @[primitives.scala 121:54]
  wire  _T_76; // @[primitives.scala 121:54]
  wire  _T_78; // @[primitives.scala 121:54]
  wire  _T_80; // @[primitives.scala 121:54]
  wire  _T_82; // @[primitives.scala 121:54]
  wire  _T_84; // @[primitives.scala 121:54]
  wire  _T_86; // @[primitives.scala 124:57]
  wire [6:0] _T_92; // @[primitives.scala 125:20]
  wire [32:0] _T_94; // @[primitives.scala 77:58]
  wire [5:0] _T_110; // @[Cat.scala 29:58]
  wire [6:0] _GEN_1; // @[MulAddRecFN.scala 125:68]
  wire [6:0] _T_111; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _T_114; // @[MulAddRecFN.scala 137:39]
  wire  _T_116; // @[MulAddRecFN.scala 137:44]
  wire  _T_118; // @[MulAddRecFN.scala 138:39]
  wire  _T_119; // @[MulAddRecFN.scala 138:44]
  wire  _T_120; // @[MulAddRecFN.scala 136:16]
  wire [74:0] _T_121; // @[Cat.scala 29:58]
  wire [75:0] alignedSigC; // @[Cat.scala 29:58]
  wire  _T_125; // @[common.scala 81:46]
  wire  _T_128; // @[common.scala 81:46]
  wire  _T_129; // @[MulAddRecFN.scala 149:32]
  wire  _T_132; // @[common.scala 81:46]
  wire [10:0] _T_137; // @[MulAddRecFN.scala 161:53]
  wire [10:0] _T_138; // @[MulAddRecFN.scala 161:12]
  assign rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[22:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[22:0]}; // @[Cat.scala 29:58]
  assign rawC_isZero = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_36 = io_c[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC_isNaN = _T_36 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC_sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC_sExp = {1'b0,$signed(io_c[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_sig = {1'h0,~rawC_isZero,io_c[22:0]}; // @[Cat.scala 29:58]
  assign signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_T_50) - 11'she5; // @[MulAddRecFN.scala 101:32]
  assign doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign _GEN_0 = {{1{rawC_sExp[9]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42]
  assign _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _T_58 = $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50]
  assign _T_60 = posNatCAlignDist <= 10'h18; // @[MulAddRecFN.scala 111:60]
  assign _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 111:23]
  assign _T_62 = posNatCAlignDist < 10'h4a; // @[MulAddRecFN.scala 115:34]
  assign _T_64 = _T_62 ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 7'h0 : _T_64; // @[MulAddRecFN.scala 113:12]
  assign _T_66 = doSubMags ? ~rawC_sig : rawC_sig; // @[MulAddRecFN.scala 121:16]
  assign _T_68 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 71:12]
  assign _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _T_71 = {rawC_sig, 2'h0}; // @[MulAddRecFN.scala 125:30]
  assign _T_74 = _T_71[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_76 = _T_71[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_78 = _T_71[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_80 = _T_71[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_82 = _T_71[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_84 = _T_71[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_86 = _T_71[26:24] != 3'h0; // @[primitives.scala 124:57]
  assign _T_92 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76,_T_74}; // @[primitives.scala 125:20]
  assign _T_94 = -33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 77:58]
  assign _T_110 = {_T_94[14],_T_94[15],_T_94[16],_T_94[17],_T_94[18],_T_94[19]}; // @[Cat.scala 29:58]
  assign _GEN_1 = {{1'd0}, _T_110}; // @[MulAddRecFN.scala 125:68]
  assign _T_111 = _T_92 & _GEN_1; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = _T_111 != 7'h0; // @[MulAddRecFN.scala 133:11]
  assign _T_114 = mainAlignedSigC[2:0] == 3'h7; // @[MulAddRecFN.scala 137:39]
  assign _T_116 = _T_114 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _T_118 = mainAlignedSigC[2:0] != 3'h0; // @[MulAddRecFN.scala 138:39]
  assign _T_119 = _T_118 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign _T_120 = doSubMags ? _T_116 : _T_119; // @[MulAddRecFN.scala 136:16]
  assign _T_121 = mainAlignedSigC[77:3]; // @[Cat.scala 29:58]
  assign alignedSigC = {_T_121,_T_120}; // @[Cat.scala 29:58]
  assign _T_125 = rawA_isNaN & ~rawA_sig[22]; // @[common.scala 81:46]
  assign _T_128 = rawB_isNaN & ~rawB_sig[22]; // @[common.scala 81:46]
  assign _T_129 = _T_125 | _T_128; // @[MulAddRecFN.scala 149:32]
  assign _T_132 = rawC_isNaN & ~rawC_sig[22]; // @[common.scala 81:46]
  assign _T_137 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53]
  assign _T_138 = CIsDominant ? $signed({{1{rawC_sExp[9]}},rawC_sExp}) : $signed(_T_137); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[23:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[23:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_129 | _T_132; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_4 & ~io_a[29]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[31:29] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_20 & ~io_b[29]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[31:29] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_36 & io_c[29]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_36 & ~io_c[29]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[31:29] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_138[9:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [9:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [4:0]  io_fromPreMul_CDom_CAlignDist,
  input  [25:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [48:0] io_mulAddResult,
  input  [2:0]  io_roundingMode,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [25:0] _T_2; // @[MulAddRecFN.scala 195:47]
  wire [25:0] _T_3; // @[MulAddRecFN.scala 194:16]
  wire [74:0] sigSum; // @[Cat.scala 29:58]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69]
  wire [9:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [9:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [49:0] _T_14; // @[Cat.scala 29:58]
  wire [49:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _T_17; // @[MulAddRecFN.scala 217:36]
  wire  _T_19; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [80:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [80:0] _T_20; // @[MulAddRecFN.scala 221:24]
  wire [28:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [26:0] _T_22; // @[MulAddRecFN.scala 224:53]
  wire  _T_25; // @[primitives.scala 121:54]
  wire  _T_27; // @[primitives.scala 121:54]
  wire  _T_29; // @[primitives.scala 121:54]
  wire  _T_31; // @[primitives.scala 121:54]
  wire  _T_33; // @[primitives.scala 121:54]
  wire  _T_35; // @[primitives.scala 121:54]
  wire  _T_37; // @[primitives.scala 124:57]
  wire [6:0] _T_43; // @[primitives.scala 125:20]
  wire [8:0] _T_46; // @[primitives.scala 77:58]
  wire [5:0] _T_62; // @[Cat.scala 29:58]
  wire [6:0] _GEN_2; // @[MulAddRecFN.scala 224:72]
  wire [6:0] _T_63; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire  _T_66; // @[MulAddRecFN.scala 228:32]
  wire  _T_67; // @[MulAddRecFN.scala 228:36]
  wire  _T_68; // @[MulAddRecFN.scala 228:61]
  wire [26:0] CDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [50:0] _GEN_3; // @[MulAddRecFN.scala 238:41]
  wire [50:0] _T_73; // @[MulAddRecFN.scala 238:41]
  wire [50:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  _T_76; // @[primitives.scala 104:54]
  wire  _T_78; // @[primitives.scala 104:54]
  wire  _T_80; // @[primitives.scala 104:54]
  wire  _T_82; // @[primitives.scala 104:54]
  wire  _T_84; // @[primitives.scala 104:54]
  wire  _T_86; // @[primitives.scala 104:54]
  wire  _T_88; // @[primitives.scala 104:54]
  wire  _T_90; // @[primitives.scala 104:54]
  wire  _T_92; // @[primitives.scala 104:54]
  wire  _T_94; // @[primitives.scala 104:54]
  wire  _T_96; // @[primitives.scala 104:54]
  wire  _T_98; // @[primitives.scala 104:54]
  wire  _T_100; // @[primitives.scala 104:54]
  wire  _T_102; // @[primitives.scala 104:54]
  wire  _T_104; // @[primitives.scala 104:54]
  wire  _T_106; // @[primitives.scala 104:54]
  wire  _T_108; // @[primitives.scala 104:54]
  wire  _T_110; // @[primitives.scala 104:54]
  wire  _T_112; // @[primitives.scala 104:54]
  wire  _T_114; // @[primitives.scala 104:54]
  wire  _T_116; // @[primitives.scala 104:54]
  wire  _T_118; // @[primitives.scala 104:54]
  wire  _T_120; // @[primitives.scala 104:54]
  wire  _T_122; // @[primitives.scala 104:54]
  wire  _T_124; // @[primitives.scala 104:54]
  wire [5:0] _T_131; // @[primitives.scala 108:20]
  wire [12:0] _T_138; // @[primitives.scala 108:20]
  wire [5:0] _T_143; // @[primitives.scala 108:20]
  wire [25:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [4:0] _T_177; // @[Mux.scala 47:69]
  wire [4:0] _T_178; // @[Mux.scala 47:69]
  wire [4:0] _T_179; // @[Mux.scala 47:69]
  wire [4:0] _T_180; // @[Mux.scala 47:69]
  wire [4:0] _T_181; // @[Mux.scala 47:69]
  wire [4:0] _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_187; // @[Mux.scala 47:69]
  wire [4:0] _T_188; // @[Mux.scala 47:69]
  wire [4:0] _T_189; // @[Mux.scala 47:69]
  wire [4:0] _T_190; // @[Mux.scala 47:69]
  wire [4:0] _T_191; // @[Mux.scala 47:69]
  wire [4:0] _T_192; // @[Mux.scala 47:69]
  wire [4:0] _T_193; // @[Mux.scala 47:69]
  wire [4:0] _T_194; // @[Mux.scala 47:69]
  wire [4:0] _T_195; // @[Mux.scala 47:69]
  wire [4:0] _T_196; // @[Mux.scala 47:69]
  wire [4:0] _T_197; // @[Mux.scala 47:69]
  wire [4:0] _T_198; // @[Mux.scala 47:69]
  wire [4:0] _T_199; // @[Mux.scala 47:69]
  wire [4:0] _T_200; // @[Mux.scala 47:69]
  wire [4:0] notCDom_normDistReduced2; // @[Mux.scala 47:69]
  wire [5:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [6:0] _T_201; // @[MulAddRecFN.scala 243:69]
  wire [9:0] _GEN_4; // @[MulAddRecFN.scala 243:46]
  wire [9:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [113:0] _GEN_5; // @[MulAddRecFN.scala 245:27]
  wire [113:0] _T_204; // @[MulAddRecFN.scala 245:27]
  wire [28:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  _T_209; // @[primitives.scala 104:54]
  wire  _T_211; // @[primitives.scala 104:54]
  wire  _T_213; // @[primitives.scala 104:54]
  wire  _T_215; // @[primitives.scala 104:54]
  wire  _T_217; // @[primitives.scala 104:54]
  wire  _T_219; // @[primitives.scala 104:54]
  wire [6:0] _T_227; // @[primitives.scala 108:20]
  wire [16:0] _T_230; // @[primitives.scala 77:58]
  wire [5:0] _T_246; // @[Cat.scala 29:58]
  wire [6:0] _GEN_6; // @[MulAddRecFN.scala 249:78]
  wire [6:0] _T_247; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire  _T_250; // @[MulAddRecFN.scala 254:35]
  wire  _T_251; // @[MulAddRecFN.scala 254:39]
  wire [26:0] notCDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _T_253; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _T_254; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _T_255; // @[MulAddRecFN.scala 274:31]
  wire  _T_256; // @[MulAddRecFN.scala 273:35]
  wire  _T_257; // @[MulAddRecFN.scala 275:32]
  wire  _T_258; // @[MulAddRecFN.scala 274:57]
  wire  _T_261; // @[MulAddRecFN.scala 276:36]
  wire  _T_262; // @[MulAddRecFN.scala 277:61]
  wire  _T_263; // @[MulAddRecFN.scala 278:35]
  wire  _T_267; // @[MulAddRecFN.scala 285:42]
  wire  _T_269; // @[MulAddRecFN.scala 287:27]
  wire  _T_270; // @[MulAddRecFN.scala 288:31]
  wire  _T_271; // @[MulAddRecFN.scala 287:54]
  wire  _T_273; // @[MulAddRecFN.scala 289:26]
  wire  _T_274; // @[MulAddRecFN.scala 289:48]
  wire  _T_275; // @[MulAddRecFN.scala 290:36]
  wire  _T_276; // @[MulAddRecFN.scala 288:43]
  wire  _T_277; // @[MulAddRecFN.scala 291:26]
  wire  _T_278; // @[MulAddRecFN.scala 292:37]
  wire  _T_279; // @[MulAddRecFN.scala 291:46]
  wire  _T_280; // @[MulAddRecFN.scala 290:48]
  wire  _T_283; // @[MulAddRecFN.scala 293:28]
  wire  _T_284; // @[MulAddRecFN.scala 294:17]
  wire  _T_285; // @[MulAddRecFN.scala 293:49]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47]
  assign _T_3 = io_mulAddResult[48] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum = {_T_3,io_mulAddResult[47:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{8{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[25:24],sigSum[72:26]}; // @[Cat.scala 29:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[74:25] : _T_14; // @[MulAddRecFN.scala 207:12]
  assign _T_17 = ~sigSum[24:1] != 24'h0; // @[MulAddRecFN.scala 217:36]
  assign _T_19 = sigSum[25:1] != 25'h0; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _T_20[49:21]; // @[MulAddRecFN.scala 221:56]
  assign _T_22 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53]
  assign _T_25 = _T_22[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_27 = _T_22[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_29 = _T_22[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_31 = _T_22[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_33 = _T_22[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_35 = _T_22[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_37 = _T_22[26:24] != 3'h0; // @[primitives.scala 124:57]
  assign _T_43 = {_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25}; // @[primitives.scala 125:20]
  assign _T_46 = -9'sh100 >>> ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 77:58]
  assign _T_62 = {_T_46[1],_T_46[2],_T_46[3],_T_46[4],_T_46[5],_T_46[6]}; // @[Cat.scala 29:58]
  assign _GEN_2 = {{1'd0}, _T_62}; // @[MulAddRecFN.scala 224:72]
  assign _T_63 = _T_43 & _GEN_2; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = _T_63 != 7'h0; // @[MulAddRecFN.scala 225:73]
  assign _T_66 = CDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 228:32]
  assign _T_67 = _T_66 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign _T_68 = _T_67 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_mainSig[28:3],_T_68}; // @[Cat.scala 29:58]
  assign notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _T_73 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[50:0] : _T_73; // @[MulAddRecFN.scala 236:12]
  assign _T_76 = notCDom_absSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_78 = notCDom_absSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_80 = notCDom_absSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_82 = notCDom_absSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_84 = notCDom_absSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_86 = notCDom_absSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_88 = notCDom_absSigSum[13:12] != 2'h0; // @[primitives.scala 104:54]
  assign _T_90 = notCDom_absSigSum[15:14] != 2'h0; // @[primitives.scala 104:54]
  assign _T_92 = notCDom_absSigSum[17:16] != 2'h0; // @[primitives.scala 104:54]
  assign _T_94 = notCDom_absSigSum[19:18] != 2'h0; // @[primitives.scala 104:54]
  assign _T_96 = notCDom_absSigSum[21:20] != 2'h0; // @[primitives.scala 104:54]
  assign _T_98 = notCDom_absSigSum[23:22] != 2'h0; // @[primitives.scala 104:54]
  assign _T_100 = notCDom_absSigSum[25:24] != 2'h0; // @[primitives.scala 104:54]
  assign _T_102 = notCDom_absSigSum[27:26] != 2'h0; // @[primitives.scala 104:54]
  assign _T_104 = notCDom_absSigSum[29:28] != 2'h0; // @[primitives.scala 104:54]
  assign _T_106 = notCDom_absSigSum[31:30] != 2'h0; // @[primitives.scala 104:54]
  assign _T_108 = notCDom_absSigSum[33:32] != 2'h0; // @[primitives.scala 104:54]
  assign _T_110 = notCDom_absSigSum[35:34] != 2'h0; // @[primitives.scala 104:54]
  assign _T_112 = notCDom_absSigSum[37:36] != 2'h0; // @[primitives.scala 104:54]
  assign _T_114 = notCDom_absSigSum[39:38] != 2'h0; // @[primitives.scala 104:54]
  assign _T_116 = notCDom_absSigSum[41:40] != 2'h0; // @[primitives.scala 104:54]
  assign _T_118 = notCDom_absSigSum[43:42] != 2'h0; // @[primitives.scala 104:54]
  assign _T_120 = notCDom_absSigSum[45:44] != 2'h0; // @[primitives.scala 104:54]
  assign _T_122 = notCDom_absSigSum[47:46] != 2'h0; // @[primitives.scala 104:54]
  assign _T_124 = notCDom_absSigSum[49:48] != 2'h0; // @[primitives.scala 104:54]
  assign _T_131 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76}; // @[primitives.scala 108:20]
  assign _T_138 = {_T_100,_T_98,_T_96,_T_94,_T_92,_T_90,_T_88,_T_131}; // @[primitives.scala 108:20]
  assign _T_143 = {_T_112,_T_110,_T_108,_T_106,_T_104,_T_102}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {notCDom_absSigSum[50],_T_124,_T_122,_T_120,_T_118,_T_116,_T_114,_T_143,_T_138}; // @[primitives.scala 108:20]
  assign _T_177 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[Mux.scala 47:69]
  assign _T_178 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _T_177; // @[Mux.scala 47:69]
  assign _T_179 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _T_178; // @[Mux.scala 47:69]
  assign _T_180 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _T_179; // @[Mux.scala 47:69]
  assign _T_181 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _T_180; // @[Mux.scala 47:69]
  assign _T_182 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _T_181; // @[Mux.scala 47:69]
  assign _T_183 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _T_182; // @[Mux.scala 47:69]
  assign _T_184 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _T_183; // @[Mux.scala 47:69]
  assign _T_185 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _T_184; // @[Mux.scala 47:69]
  assign _T_186 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _T_185; // @[Mux.scala 47:69]
  assign _T_187 = notCDom_reduced2AbsSigSum[11] ? 5'he : _T_186; // @[Mux.scala 47:69]
  assign _T_188 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _T_187; // @[Mux.scala 47:69]
  assign _T_189 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _T_188; // @[Mux.scala 47:69]
  assign _T_190 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _T_189; // @[Mux.scala 47:69]
  assign _T_191 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _T_190; // @[Mux.scala 47:69]
  assign _T_192 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _T_191; // @[Mux.scala 47:69]
  assign _T_193 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _T_192; // @[Mux.scala 47:69]
  assign _T_194 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _T_193; // @[Mux.scala 47:69]
  assign _T_195 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _T_194; // @[Mux.scala 47:69]
  assign _T_196 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _T_195; // @[Mux.scala 47:69]
  assign _T_197 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _T_196; // @[Mux.scala 47:69]
  assign _T_198 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _T_197; // @[Mux.scala 47:69]
  assign _T_199 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _T_198; // @[Mux.scala 47:69]
  assign _T_200 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _T_199; // @[Mux.scala 47:69]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _T_200; // @[Mux.scala 47:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _T_201 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_4 = {{3{_T_201[6]}},_T_201}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46]
  assign _GEN_5 = {{63'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _T_204 = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _T_204[51:23]; // @[MulAddRecFN.scala 245:50]
  assign _T_209 = notCDom_reduced2AbsSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_211 = notCDom_reduced2AbsSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_213 = notCDom_reduced2AbsSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_215 = notCDom_reduced2AbsSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_217 = notCDom_reduced2AbsSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_219 = notCDom_reduced2AbsSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_227 = {notCDom_reduced2AbsSigSum[12],_T_219,_T_217,_T_215,_T_213,_T_211,_T_209}; // @[primitives.scala 108:20]
  assign _T_230 = -17'sh10000 >>> ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 77:58]
  assign _T_246 = {_T_230[1],_T_230[2],_T_230[3],_T_230[4],_T_230[5],_T_230[6]}; // @[Cat.scala 29:58]
  assign _GEN_6 = {{1'd0}, _T_246}; // @[MulAddRecFN.scala 249:78]
  assign _T_247 = _T_227 & _GEN_6; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = _T_247 != 7'h0; // @[MulAddRecFN.scala 251:11]
  assign _T_250 = notCDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 254:35]
  assign _T_251 = _T_250 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_mainSig[28:3],_T_251}; // @[Cat.scala 29:58]
  assign notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _T_253 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_253; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _T_254 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _T_254 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _T_255 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _T_256 = io_fromPreMul_isSigNaNAny | _T_255; // @[MulAddRecFN.scala 273:35]
  assign _T_257 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _T_258 = _T_256 | _T_257; // @[MulAddRecFN.scala 274:57]
  assign _T_261 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _T_262 = _T_261 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _T_263 = _T_262 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _T_267 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _T_269 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _T_270 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _T_271 = _T_269 | _T_270; // @[MulAddRecFN.scala 287:54]
  assign _T_273 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _T_274 = _T_273 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _T_275 = _T_274 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _T_276 = _T_271 | _T_275; // @[MulAddRecFN.scala 288:43]
  assign _T_277 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _T_278 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _T_279 = _T_277 & _T_278; // @[MulAddRecFN.scala 291:46]
  assign _T_280 = _T_276 | _T_279; // @[MulAddRecFN.scala 290:48]
  assign _T_283 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _T_284 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _T_285 = _T_283 & _T_284; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_258 | _T_263; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_267; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_280 | _T_285; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  _T_5; // @[primitives.scala 57:25]
  wire  _T_7; // @[primitives.scala 57:25]
  wire  _T_9; // @[primitives.scala 57:25]
  wire [5:0] _T_10; // @[primitives.scala 58:26]
  wire [64:0] _T_11; // @[primitives.scala 77:58]
  wire [15:0] _T_17; // @[Bitwise.scala 102:31]
  wire [15:0] _T_19; // @[Bitwise.scala 102:65]
  wire [15:0] _T_21; // @[Bitwise.scala 102:75]
  wire [15:0] _T_22; // @[Bitwise.scala 102:39]
  wire [15:0] _GEN_0; // @[Bitwise.scala 102:31]
  wire [15:0] _T_27; // @[Bitwise.scala 102:31]
  wire [15:0] _T_29; // @[Bitwise.scala 102:65]
  wire [15:0] _T_31; // @[Bitwise.scala 102:75]
  wire [15:0] _T_32; // @[Bitwise.scala 102:39]
  wire [15:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [15:0] _T_37; // @[Bitwise.scala 102:31]
  wire [15:0] _T_39; // @[Bitwise.scala 102:65]
  wire [15:0] _T_41; // @[Bitwise.scala 102:75]
  wire [15:0] _T_42; // @[Bitwise.scala 102:39]
  wire [15:0] _GEN_2; // @[Bitwise.scala 102:31]
  wire [15:0] _T_47; // @[Bitwise.scala 102:31]
  wire [15:0] _T_49; // @[Bitwise.scala 102:65]
  wire [15:0] _T_51; // @[Bitwise.scala 102:75]
  wire [15:0] _T_52; // @[Bitwise.scala 102:39]
  wire [21:0] _T_69; // @[Cat.scala 29:58]
  wire [21:0] _T_71; // @[primitives.scala 74:21]
  wire [24:0] _T_73; // @[Cat.scala 29:58]
  wire [2:0] _T_83; // @[Cat.scala 29:58]
  wire [2:0] _T_84; // @[primitives.scala 61:24]
  wire [24:0] _T_85; // @[primitives.scala 66:24]
  wire [24:0] _T_86; // @[primitives.scala 61:24]
  wire [24:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [24:0] _T_87; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [26:0] _T_88; // @[Cat.scala 29:58]
  wire [26:0] _T_90; // @[Cat.scala 29:58]
  wire [26:0] _T_92; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _T_93; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_94; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _T_95; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_96; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_97; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_98; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_99; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_100; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_101; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _T_102; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _T_104; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_105; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_107; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _T_109; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _T_111; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _T_113; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_115; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _T_117; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_118; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _T_119; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_121; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_5; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] _T_122; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_127; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_132; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _T_134; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _T_136; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_137; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _T_139; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_140; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_141; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  _T_144; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _T_145; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_146; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_147; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_150; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _T_151; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_155; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _T_157; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_158; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_159; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_160; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_162; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _T_167; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_169; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_171; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_175; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _T_176; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _T_178; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _T_180; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _T_182; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _T_183; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _T_185; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _T_189; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _T_190; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _T_191; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _T_192; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _T_193; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _T_194; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _T_195; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_196; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_197; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _T_198; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _T_199; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _T_201; // @[Bitwise.scala 71:12]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] _T_202; // @[Cat.scala 29:58]
  wire [1:0] _T_204; // @[Cat.scala 29:58]
  wire [2:0] _T_206; // @[Cat.scala 29:58]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign _T_5 = ~io_in_sExp[8]; // @[primitives.scala 57:25]
  assign _T_7 = ~io_in_sExp[7]; // @[primitives.scala 57:25]
  assign _T_9 = ~io_in_sExp[6]; // @[primitives.scala 57:25]
  assign _T_10 = ~io_in_sExp[5:0]; // @[primitives.scala 58:26]
  assign _T_11 = -65'sh10000000000000000 >>> _T_10; // @[primitives.scala 77:58]
  assign _T_17 = {{8'd0}, _T_11[57:50]}; // @[Bitwise.scala 102:31]
  assign _T_19 = {_T_11[49:42], 8'h0}; // @[Bitwise.scala 102:65]
  assign _T_21 = _T_19 & 16'hff00; // @[Bitwise.scala 102:75]
  assign _T_22 = _T_17 | _T_21; // @[Bitwise.scala 102:39]
  assign _GEN_0 = {{4'd0}, _T_22[15:4]}; // @[Bitwise.scala 102:31]
  assign _T_27 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 102:31]
  assign _T_29 = {_T_22[11:0], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_31 = _T_29 & 16'hf0f0; // @[Bitwise.scala 102:75]
  assign _T_32 = _T_27 | _T_31; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{2'd0}, _T_32[15:2]}; // @[Bitwise.scala 102:31]
  assign _T_37 = _GEN_1 & 16'h3333; // @[Bitwise.scala 102:31]
  assign _T_39 = {_T_32[13:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_41 = _T_39 & 16'hcccc; // @[Bitwise.scala 102:75]
  assign _T_42 = _T_37 | _T_41; // @[Bitwise.scala 102:39]
  assign _GEN_2 = {{1'd0}, _T_42[15:1]}; // @[Bitwise.scala 102:31]
  assign _T_47 = _GEN_2 & 16'h5555; // @[Bitwise.scala 102:31]
  assign _T_49 = {_T_42[14:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_51 = _T_49 & 16'haaaa; // @[Bitwise.scala 102:75]
  assign _T_52 = _T_47 | _T_51; // @[Bitwise.scala 102:39]
  assign _T_69 = {_T_52,_T_11[58],_T_11[59],_T_11[60],_T_11[61],_T_11[62],_T_11[63]}; // @[Cat.scala 29:58]
  assign _T_71 = _T_9 ? 22'h0 : ~_T_69; // @[primitives.scala 74:21]
  assign _T_73 = {~_T_71,3'h7}; // @[Cat.scala 29:58]
  assign _T_83 = {_T_11[0],_T_11[1],_T_11[2]}; // @[Cat.scala 29:58]
  assign _T_84 = _T_9 ? _T_83 : 3'h0; // @[primitives.scala 61:24]
  assign _T_85 = _T_7 ? _T_73 : {{22'd0}, _T_84}; // @[primitives.scala 66:24]
  assign _T_86 = _T_5 ? _T_85 : 25'h0; // @[primitives.scala 61:24]
  assign _GEN_3 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_87 = _T_86 | _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_88 = {_T_87,2'h3}; // @[Cat.scala 29:58]
  assign _T_90 = {1'h0,_T_88[26:1]}; // @[Cat.scala 29:58]
  assign _T_92 = ~_T_90 & _T_88; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_93 = io_in_sig & _T_92; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_94 = _T_93 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_95 = io_in_sig & _T_90; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_96 = _T_95 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_97 = _T_94 | _T_96; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_98 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_99 = _T_98 & _T_94; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_100 = roundMagUp & _T_97; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_101 = _T_99 | _T_100; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_102 = io_in_sig | _T_88; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_104 = _T_102[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_105 = roundingMode_near_even & _T_94; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_107 = _T_105 & ~_T_96; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_109 = _T_107 ? _T_88[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_111 = _T_104 & ~_T_109; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_113 = io_in_sig & ~_T_88; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_115 = roundingMode_odd & _T_97; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_117 = _T_115 ? _T_92[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_4 = {{1'd0}, _T_113[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_118 = _GEN_4 | _T_117; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_119 = _T_101 ? _T_111 : _T_118; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_121 = {1'b0,$signed(_T_119[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_5 = {{7{_T_121[2]}},_T_121}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_122 = $signed(io_in_sExp) + $signed(_GEN_5); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_122[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? _T_119[23:1] : _T_119[22:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _T_127 = _T_122[10:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_127) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_122) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_132 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _T_134 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _T_136 = io_in_sig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_137 = _T_134 | _T_136; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _T_139 = _T_98 & _T_132; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_140 = roundMagUp & _T_137; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_141 = _T_139 | _T_140; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_144 = doShiftSigDown1 ? _T_119[25] : _T_119[24]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _T_145 = io_in_sExp[9:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_146 = $signed(_T_145) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_147 = _T_97 & _T_146; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_150 = doShiftSigDown1 ? _T_88[3] : _T_88[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _T_151 = _T_147 & _T_150; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_155 = doShiftSigDown1 ? _T_88[4] : _T_88[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _T_157 = io_detectTininess & ~_T_155; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_158 = _T_157 & _T_144; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_159 = _T_158 & _T_94; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_160 = _T_159 & _T_141; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_162 = _T_151 & ~_T_160; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_162; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_97; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign _T_167 = ~isNaNOut & ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_167 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_169 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_169; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_98 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_171 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_172 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_171 & _T_172; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_174 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = io_in_isInf | _T_174; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_175 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_176 = _T_175 ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_178 = common_expOut & ~_T_176; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_180 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_182 = _T_178 & ~_T_180; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_183 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_185 = _T_182 & ~_T_183; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_186 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_188 = _T_185 & ~_T_186; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_189 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_190 = _T_188 | _T_189; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_191 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_192 = _T_190 | _T_191; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_193 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_194 = _T_192 | _T_193; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_195 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_194 | _T_195; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_196 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_197 = _T_196 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_198 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_199 = _T_197 ? _T_198 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_201 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 71:12]
  assign fractOut = _T_199 | _T_201; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_202 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_204 = {underflow,inexact}; // @[Cat.scala 29:58]
  assign _T_206 = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_202,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_206,_T_204}; // @[RoundAnyRawFNToRecFN.scala 285:23]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
endmodule
module MulAddRecFN(
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[MulAddRecFN.scala 318:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[MulAddRecFN.scala 318:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[MulAddRecFN.scala 318:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[MulAddRecFN.scala 318:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 318:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 318:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 318:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 318:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 320:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 320:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 320:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[MulAddRecFN.scala 320:15]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 320:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 320:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 320:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulAddRecFN.scala 340:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[MulAddRecFN.scala 340:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[MulAddRecFN.scala 340:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[MulAddRecFN.scala 340:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 340:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[MulAddRecFN.scala 340:15]
  wire [47:0] _T; // @[MulAddRecFN.scala 328:45]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[MulAddRecFN.scala 318:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[MulAddRecFN.scala 320:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[MulAddRecFN.scala 340:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags)
  );
  assign _T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 328:45]
  assign io_out = roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 346:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[MulAddRecFN.scala 347:23]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[MulAddRecFN.scala 323:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[MulAddRecFN.scala 324:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[MulAddRecFN.scala 325:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 334:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = io_roundingMode; // @[MulAddRecFN.scala 335:46]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 341:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_roundingMode = io_roundingMode; // @[MulAddRecFN.scala 344:39]
  assign roundRawFNToRecFN_io_detectTininess = io_detectTininess; // @[MulAddRecFN.scala 345:41]
endmodule
module ValExec_MulAddRecF32(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  input  [31:0] io_c,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [31:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [32:0] io_expected_recOut,
  output [32:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [32:0] mulAddRecFN_io_a; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [32:0] mulAddRecFN_io_b; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [32:0] mulAddRecFN_io_c; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [2:0] mulAddRecFN_io_roundingMode; // @[ValExec_MulAddRecFN.scala 66:29]
  wire  mulAddRecFN_io_detectTininess; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [32:0] mulAddRecFN_io_out; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [4:0] mulAddRecFN_io_exceptionFlags; // @[ValExec_MulAddRecFN.scala 66:29]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_48; // @[Mux.scala 47:69]
  wire [4:0] _T_49; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61; // @[rawFloatFromFN.scala 63:62]
  wire  _T_64; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_67; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_69; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_71; // @[Cat.scala 29:58]
  wire [2:0] _T_73; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_75; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_78; // @[Cat.scala 29:58]
  wire [3:0] _T_79; // @[Cat.scala 29:58]
  wire  _T_84; // @[rawFloatFromFN.scala 50:34]
  wire  _T_85; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_120; // @[Mux.scala 47:69]
  wire [4:0] _T_121; // @[Mux.scala 47:69]
  wire [4:0] _T_122; // @[Mux.scala 47:69]
  wire [4:0] _T_123; // @[Mux.scala 47:69]
  wire [4:0] _T_124; // @[Mux.scala 47:69]
  wire [4:0] _T_125; // @[Mux.scala 47:69]
  wire [4:0] _T_126; // @[Mux.scala 47:69]
  wire [4:0] _T_127; // @[Mux.scala 47:69]
  wire [4:0] _T_128; // @[Mux.scala 47:69]
  wire [4:0] _T_129; // @[Mux.scala 47:69]
  wire [4:0] _T_130; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_131; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_133; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_134; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_135; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_136; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_137; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_139; // @[rawFloatFromFN.scala 59:15]
  wire  _T_140; // @[rawFloatFromFN.scala 62:34]
  wire  _T_142; // @[rawFloatFromFN.scala 63:62]
  wire  _T_145; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_148; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_150; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_152; // @[Cat.scala 29:58]
  wire [2:0] _T_154; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_156; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_159; // @[Cat.scala 29:58]
  wire [3:0] _T_160; // @[Cat.scala 29:58]
  wire  _T_165; // @[rawFloatFromFN.scala 50:34]
  wire  _T_166; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_190; // @[Mux.scala 47:69]
  wire [4:0] _T_191; // @[Mux.scala 47:69]
  wire [4:0] _T_192; // @[Mux.scala 47:69]
  wire [4:0] _T_193; // @[Mux.scala 47:69]
  wire [4:0] _T_194; // @[Mux.scala 47:69]
  wire [4:0] _T_195; // @[Mux.scala 47:69]
  wire [4:0] _T_196; // @[Mux.scala 47:69]
  wire [4:0] _T_197; // @[Mux.scala 47:69]
  wire [4:0] _T_198; // @[Mux.scala 47:69]
  wire [4:0] _T_199; // @[Mux.scala 47:69]
  wire [4:0] _T_200; // @[Mux.scala 47:69]
  wire [4:0] _T_201; // @[Mux.scala 47:69]
  wire [4:0] _T_202; // @[Mux.scala 47:69]
  wire [4:0] _T_203; // @[Mux.scala 47:69]
  wire [4:0] _T_204; // @[Mux.scala 47:69]
  wire [4:0] _T_205; // @[Mux.scala 47:69]
  wire [4:0] _T_206; // @[Mux.scala 47:69]
  wire [4:0] _T_207; // @[Mux.scala 47:69]
  wire [4:0] _T_208; // @[Mux.scala 47:69]
  wire [4:0] _T_209; // @[Mux.scala 47:69]
  wire [4:0] _T_210; // @[Mux.scala 47:69]
  wire [4:0] _T_211; // @[Mux.scala 47:69]
  wire [53:0] _GEN_10; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_212; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_214; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_11; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_215; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_216; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_217; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_12; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_218; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_13; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_220; // @[rawFloatFromFN.scala 59:15]
  wire  _T_221; // @[rawFloatFromFN.scala 62:34]
  wire  _T_223; // @[rawFloatFromFN.scala 63:62]
  wire  _T_226; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_229; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_231; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_233; // @[Cat.scala 29:58]
  wire [2:0] _T_235; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_14; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_237; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_240; // @[Cat.scala 29:58]
  wire [3:0] _T_241; // @[Cat.scala 29:58]
  wire  _T_246; // @[rawFloatFromFN.scala 50:34]
  wire  _T_247; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_271; // @[Mux.scala 47:69]
  wire [4:0] _T_272; // @[Mux.scala 47:69]
  wire [4:0] _T_273; // @[Mux.scala 47:69]
  wire [4:0] _T_274; // @[Mux.scala 47:69]
  wire [4:0] _T_275; // @[Mux.scala 47:69]
  wire [4:0] _T_276; // @[Mux.scala 47:69]
  wire [4:0] _T_277; // @[Mux.scala 47:69]
  wire [4:0] _T_278; // @[Mux.scala 47:69]
  wire [4:0] _T_279; // @[Mux.scala 47:69]
  wire [4:0] _T_280; // @[Mux.scala 47:69]
  wire [4:0] _T_281; // @[Mux.scala 47:69]
  wire [4:0] _T_282; // @[Mux.scala 47:69]
  wire [4:0] _T_283; // @[Mux.scala 47:69]
  wire [4:0] _T_284; // @[Mux.scala 47:69]
  wire [4:0] _T_285; // @[Mux.scala 47:69]
  wire [4:0] _T_286; // @[Mux.scala 47:69]
  wire [4:0] _T_287; // @[Mux.scala 47:69]
  wire [4:0] _T_288; // @[Mux.scala 47:69]
  wire [4:0] _T_289; // @[Mux.scala 47:69]
  wire [4:0] _T_290; // @[Mux.scala 47:69]
  wire [4:0] _T_291; // @[Mux.scala 47:69]
  wire [4:0] _T_292; // @[Mux.scala 47:69]
  wire [53:0] _GEN_15; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_293; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_295; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_16; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_296; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_297; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_298; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_17; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_299; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_18; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_301; // @[rawFloatFromFN.scala 59:15]
  wire  _T_302; // @[rawFloatFromFN.scala 62:34]
  wire  _T_304; // @[rawFloatFromFN.scala 63:62]
  wire  _T_307; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_310; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_312; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_314; // @[Cat.scala 29:58]
  wire [2:0] _T_316; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_19; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_318; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_321; // @[Cat.scala 29:58]
  wire [3:0] _T_322; // @[Cat.scala 29:58]
  wire  _T_327; // @[tests.scala 48:26]
  wire  _T_329; // @[tests.scala 48:55]
  wire  _T_330; // @[tests.scala 48:39]
  wire  _T_331; // @[tests.scala 49:20]
  wire  _T_334; // @[tests.scala 49:54]
  wire  _T_335; // @[tests.scala 49:31]
  wire  _T_337; // @[tests.scala 50:30]
  wire  _T_339; // @[tests.scala 50:66]
  wire  _T_340; // @[tests.scala 50:16]
  wire  _T_341; // @[tests.scala 48:12]
  wire  _T_342; // @[ValExec_MulAddRecFN.scala 82:35]
  MulAddRecFN mulAddRecFN ( // @[ValExec_MulAddRecFN.scala 66:29]
    .io_a(mulAddRecFN_io_a),
    .io_b(mulAddRecFN_io_b),
    .io_c(mulAddRecFN_io_c),
    .io_roundingMode(mulAddRecFN_io_roundingMode),
    .io_detectTininess(mulAddRecFN_io_detectTininess),
    .io_out(mulAddRecFN_io_out),
    .io_exceptionFlags(mulAddRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  assign _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  assign _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  assign _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  assign _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  assign _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  assign _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  assign _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  assign _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  assign _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  assign _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  assign _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  assign _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  assign _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  assign _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  assign _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  assign _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  assign _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  assign _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  assign _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  assign _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  assign _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  assign _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  assign _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  assign _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  assign _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_64 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_67 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_69 = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_71 = {1'h0,~_T_59,_T_69}; // @[Cat.scala 29:58]
  assign _T_73 = _T_59 ? 3'h0 : _T_67[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_64}; // @[recFNFromFN.scala 48:79]
  assign _T_75 = _T_73 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_78 = {_T_67[5:0],_T_71[22:0]}; // @[Cat.scala 29:58]
  assign _T_79 = {io_a[31],_T_75}; // @[Cat.scala 29:58]
  assign _T_84 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_85 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_109 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_110 = io_b[2] ? 5'h14 : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = io_b[3] ? 5'h13 : _T_110; // @[Mux.scala 47:69]
  assign _T_112 = io_b[4] ? 5'h12 : _T_111; // @[Mux.scala 47:69]
  assign _T_113 = io_b[5] ? 5'h11 : _T_112; // @[Mux.scala 47:69]
  assign _T_114 = io_b[6] ? 5'h10 : _T_113; // @[Mux.scala 47:69]
  assign _T_115 = io_b[7] ? 5'hf : _T_114; // @[Mux.scala 47:69]
  assign _T_116 = io_b[8] ? 5'he : _T_115; // @[Mux.scala 47:69]
  assign _T_117 = io_b[9] ? 5'hd : _T_116; // @[Mux.scala 47:69]
  assign _T_118 = io_b[10] ? 5'hc : _T_117; // @[Mux.scala 47:69]
  assign _T_119 = io_b[11] ? 5'hb : _T_118; // @[Mux.scala 47:69]
  assign _T_120 = io_b[12] ? 5'ha : _T_119; // @[Mux.scala 47:69]
  assign _T_121 = io_b[13] ? 5'h9 : _T_120; // @[Mux.scala 47:69]
  assign _T_122 = io_b[14] ? 5'h8 : _T_121; // @[Mux.scala 47:69]
  assign _T_123 = io_b[15] ? 5'h7 : _T_122; // @[Mux.scala 47:69]
  assign _T_124 = io_b[16] ? 5'h6 : _T_123; // @[Mux.scala 47:69]
  assign _T_125 = io_b[17] ? 5'h5 : _T_124; // @[Mux.scala 47:69]
  assign _T_126 = io_b[18] ? 5'h4 : _T_125; // @[Mux.scala 47:69]
  assign _T_127 = io_b[19] ? 5'h3 : _T_126; // @[Mux.scala 47:69]
  assign _T_128 = io_b[20] ? 5'h2 : _T_127; // @[Mux.scala 47:69]
  assign _T_129 = io_b[21] ? 5'h1 : _T_128; // @[Mux.scala 47:69]
  assign _T_130 = io_b[22] ? 5'h0 : _T_129; // @[Mux.scala 47:69]
  assign _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_131 = _GEN_5 << _T_130; // @[rawFloatFromFN.scala 54:36]
  assign _T_133 = {_T_131[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{4'd0}, _T_130}; // @[rawFloatFromFN.scala 57:26]
  assign _T_134 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_135 = _T_84 ? _T_134 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_136 = _T_84 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{6'd0}, _T_136}; // @[rawFloatFromFN.scala 60:22]
  assign _T_137 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_137}; // @[rawFloatFromFN.scala 59:15]
  assign _T_139 = _T_135 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_140 = _T_84 & _T_85; // @[rawFloatFromFN.scala 62:34]
  assign _T_142 = _T_139[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_145 = _T_142 & ~_T_85; // @[rawFloatFromFN.scala 66:33]
  assign _T_148 = {1'b0,$signed(_T_139)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_150 = _T_84 ? _T_133 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_152 = {1'h0,~_T_140,_T_150}; // @[Cat.scala 29:58]
  assign _T_154 = _T_140 ? 3'h0 : _T_148[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_145}; // @[recFNFromFN.scala 48:79]
  assign _T_156 = _T_154 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_159 = {_T_148[5:0],_T_152[22:0]}; // @[Cat.scala 29:58]
  assign _T_160 = {io_b[31],_T_156}; // @[Cat.scala 29:58]
  assign _T_165 = io_c[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_166 = io_c[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_190 = io_c[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_191 = io_c[2] ? 5'h14 : _T_190; // @[Mux.scala 47:69]
  assign _T_192 = io_c[3] ? 5'h13 : _T_191; // @[Mux.scala 47:69]
  assign _T_193 = io_c[4] ? 5'h12 : _T_192; // @[Mux.scala 47:69]
  assign _T_194 = io_c[5] ? 5'h11 : _T_193; // @[Mux.scala 47:69]
  assign _T_195 = io_c[6] ? 5'h10 : _T_194; // @[Mux.scala 47:69]
  assign _T_196 = io_c[7] ? 5'hf : _T_195; // @[Mux.scala 47:69]
  assign _T_197 = io_c[8] ? 5'he : _T_196; // @[Mux.scala 47:69]
  assign _T_198 = io_c[9] ? 5'hd : _T_197; // @[Mux.scala 47:69]
  assign _T_199 = io_c[10] ? 5'hc : _T_198; // @[Mux.scala 47:69]
  assign _T_200 = io_c[11] ? 5'hb : _T_199; // @[Mux.scala 47:69]
  assign _T_201 = io_c[12] ? 5'ha : _T_200; // @[Mux.scala 47:69]
  assign _T_202 = io_c[13] ? 5'h9 : _T_201; // @[Mux.scala 47:69]
  assign _T_203 = io_c[14] ? 5'h8 : _T_202; // @[Mux.scala 47:69]
  assign _T_204 = io_c[15] ? 5'h7 : _T_203; // @[Mux.scala 47:69]
  assign _T_205 = io_c[16] ? 5'h6 : _T_204; // @[Mux.scala 47:69]
  assign _T_206 = io_c[17] ? 5'h5 : _T_205; // @[Mux.scala 47:69]
  assign _T_207 = io_c[18] ? 5'h4 : _T_206; // @[Mux.scala 47:69]
  assign _T_208 = io_c[19] ? 5'h3 : _T_207; // @[Mux.scala 47:69]
  assign _T_209 = io_c[20] ? 5'h2 : _T_208; // @[Mux.scala 47:69]
  assign _T_210 = io_c[21] ? 5'h1 : _T_209; // @[Mux.scala 47:69]
  assign _T_211 = io_c[22] ? 5'h0 : _T_210; // @[Mux.scala 47:69]
  assign _GEN_10 = {{31'd0}, io_c[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_212 = _GEN_10 << _T_211; // @[rawFloatFromFN.scala 54:36]
  assign _T_214 = {_T_212[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_11 = {{4'd0}, _T_211}; // @[rawFloatFromFN.scala 57:26]
  assign _T_215 = _GEN_11 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_216 = _T_165 ? _T_215 : {{1'd0}, io_c[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_217 = _T_165 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_12 = {{6'd0}, _T_217}; // @[rawFloatFromFN.scala 60:22]
  assign _T_218 = 8'h80 | _GEN_12; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_13 = {{1'd0}, _T_218}; // @[rawFloatFromFN.scala 59:15]
  assign _T_220 = _T_216 + _GEN_13; // @[rawFloatFromFN.scala 59:15]
  assign _T_221 = _T_165 & _T_166; // @[rawFloatFromFN.scala 62:34]
  assign _T_223 = _T_220[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_226 = _T_223 & ~_T_166; // @[rawFloatFromFN.scala 66:33]
  assign _T_229 = {1'b0,$signed(_T_220)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_231 = _T_165 ? _T_214 : io_c[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_233 = {1'h0,~_T_221,_T_231}; // @[Cat.scala 29:58]
  assign _T_235 = _T_221 ? 3'h0 : _T_229[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_14 = {{2'd0}, _T_226}; // @[recFNFromFN.scala 48:79]
  assign _T_237 = _T_235 | _GEN_14; // @[recFNFromFN.scala 48:79]
  assign _T_240 = {_T_229[5:0],_T_233[22:0]}; // @[Cat.scala 29:58]
  assign _T_241 = {io_c[31],_T_237}; // @[Cat.scala 29:58]
  assign _T_246 = io_expected_out[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_247 = io_expected_out[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_271 = io_expected_out[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_272 = io_expected_out[2] ? 5'h14 : _T_271; // @[Mux.scala 47:69]
  assign _T_273 = io_expected_out[3] ? 5'h13 : _T_272; // @[Mux.scala 47:69]
  assign _T_274 = io_expected_out[4] ? 5'h12 : _T_273; // @[Mux.scala 47:69]
  assign _T_275 = io_expected_out[5] ? 5'h11 : _T_274; // @[Mux.scala 47:69]
  assign _T_276 = io_expected_out[6] ? 5'h10 : _T_275; // @[Mux.scala 47:69]
  assign _T_277 = io_expected_out[7] ? 5'hf : _T_276; // @[Mux.scala 47:69]
  assign _T_278 = io_expected_out[8] ? 5'he : _T_277; // @[Mux.scala 47:69]
  assign _T_279 = io_expected_out[9] ? 5'hd : _T_278; // @[Mux.scala 47:69]
  assign _T_280 = io_expected_out[10] ? 5'hc : _T_279; // @[Mux.scala 47:69]
  assign _T_281 = io_expected_out[11] ? 5'hb : _T_280; // @[Mux.scala 47:69]
  assign _T_282 = io_expected_out[12] ? 5'ha : _T_281; // @[Mux.scala 47:69]
  assign _T_283 = io_expected_out[13] ? 5'h9 : _T_282; // @[Mux.scala 47:69]
  assign _T_284 = io_expected_out[14] ? 5'h8 : _T_283; // @[Mux.scala 47:69]
  assign _T_285 = io_expected_out[15] ? 5'h7 : _T_284; // @[Mux.scala 47:69]
  assign _T_286 = io_expected_out[16] ? 5'h6 : _T_285; // @[Mux.scala 47:69]
  assign _T_287 = io_expected_out[17] ? 5'h5 : _T_286; // @[Mux.scala 47:69]
  assign _T_288 = io_expected_out[18] ? 5'h4 : _T_287; // @[Mux.scala 47:69]
  assign _T_289 = io_expected_out[19] ? 5'h3 : _T_288; // @[Mux.scala 47:69]
  assign _T_290 = io_expected_out[20] ? 5'h2 : _T_289; // @[Mux.scala 47:69]
  assign _T_291 = io_expected_out[21] ? 5'h1 : _T_290; // @[Mux.scala 47:69]
  assign _T_292 = io_expected_out[22] ? 5'h0 : _T_291; // @[Mux.scala 47:69]
  assign _GEN_15 = {{31'd0}, io_expected_out[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_293 = _GEN_15 << _T_292; // @[rawFloatFromFN.scala 54:36]
  assign _T_295 = {_T_293[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_16 = {{4'd0}, _T_292}; // @[rawFloatFromFN.scala 57:26]
  assign _T_296 = _GEN_16 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_297 = _T_246 ? _T_296 : {{1'd0}, io_expected_out[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_298 = _T_246 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_17 = {{6'd0}, _T_298}; // @[rawFloatFromFN.scala 60:22]
  assign _T_299 = 8'h80 | _GEN_17; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_18 = {{1'd0}, _T_299}; // @[rawFloatFromFN.scala 59:15]
  assign _T_301 = _T_297 + _GEN_18; // @[rawFloatFromFN.scala 59:15]
  assign _T_302 = _T_246 & _T_247; // @[rawFloatFromFN.scala 62:34]
  assign _T_304 = _T_301[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_307 = _T_304 & ~_T_247; // @[rawFloatFromFN.scala 66:33]
  assign _T_310 = {1'b0,$signed(_T_301)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_312 = _T_246 ? _T_295 : io_expected_out[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_314 = {1'h0,~_T_302,_T_312}; // @[Cat.scala 29:58]
  assign _T_316 = _T_302 ? 3'h0 : _T_310[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_19 = {{2'd0}, _T_307}; // @[recFNFromFN.scala 48:79]
  assign _T_318 = _T_316 | _GEN_19; // @[recFNFromFN.scala 48:79]
  assign _T_321 = {_T_310[5:0],_T_314[22:0]}; // @[Cat.scala 29:58]
  assign _T_322 = {io_expected_out[31],_T_318}; // @[Cat.scala 29:58]
  assign _T_327 = io_actual_out[31:29] == 3'h0; // @[tests.scala 48:26]
  assign _T_329 = io_actual_out[31:29] == 3'h7; // @[tests.scala 48:55]
  assign _T_330 = _T_327 | _T_329; // @[tests.scala 48:39]
  assign _T_331 = io_actual_out[32:29] == io_expected_recOut[32:29]; // @[tests.scala 49:20]
  assign _T_334 = io_actual_out[22:0] == io_expected_recOut[22:0]; // @[tests.scala 49:54]
  assign _T_335 = _T_331 & _T_334; // @[tests.scala 49:31]
  assign _T_337 = io_actual_out[31:29] == 3'h6; // @[tests.scala 50:30]
  assign _T_339 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_340 = _T_337 ? _T_331 : _T_339; // @[tests.scala 50:16]
  assign _T_341 = _T_330 ? _T_335 : _T_340; // @[tests.scala 48:12]
  assign _T_342 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_MulAddRecFN.scala 82:35]
  assign io_expected_recOut = {_T_322,_T_321}; // @[ValExec_MulAddRecFN.scala 74:24]
  assign io_actual_out = mulAddRecFN_io_out; // @[ValExec_MulAddRecFN.scala 76:19]
  assign io_actual_exceptionFlags = mulAddRecFN_io_exceptionFlags; // @[ValExec_MulAddRecFN.scala 77:30]
  assign io_check = 1'h1; // @[ValExec_MulAddRecFN.scala 79:14]
  assign io_pass = _T_341 & _T_342; // @[ValExec_MulAddRecFN.scala 80:13]
  assign mulAddRecFN_io_a = {_T_79,_T_78}; // @[ValExec_MulAddRecFN.scala 68:22]
  assign mulAddRecFN_io_b = {_T_160,_T_159}; // @[ValExec_MulAddRecFN.scala 69:22]
  assign mulAddRecFN_io_c = {_T_241,_T_240}; // @[ValExec_MulAddRecFN.scala 70:22]
  assign mulAddRecFN_io_roundingMode = io_roundingMode; // @[ValExec_MulAddRecFN.scala 71:35]
  assign mulAddRecFN_io_detectTininess = io_detectTininess; // @[ValExec_MulAddRecFN.scala 72:35]
endmodule
