module MulAddRecFNToRaw_preMul(
  input  [64:0]  io_a,
  input  [64:0]  io_b,
  input  [64:0]  io_c,
  output [52:0]  io_mulAddA,
  output [52:0]  io_mulAddB,
  output [105:0] io_mulAddC,
  output         io_toPostMul_isSigNaNAny,
  output         io_toPostMul_isNaNAOrB,
  output         io_toPostMul_isInfA,
  output         io_toPostMul_isZeroA,
  output         io_toPostMul_isInfB,
  output         io_toPostMul_isZeroB,
  output         io_toPostMul_signProd,
  output         io_toPostMul_isNaNC,
  output         io_toPostMul_isInfC,
  output         io_toPostMul_isZeroC,
  output [12:0]  io_toPostMul_sExpSum,
  output         io_toPostMul_doSubMags,
  output         io_toPostMul_CIsDominant,
  output [5:0]   io_toPostMul_CDom_CAlignDist,
  output [54:0]  io_toPostMul_highAlignedSigC,
  output         io_toPostMul_bit0AlignedSigC
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawB_sig; // @[Cat.scala 29:58]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_36; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawC_sig; // @[Cat.scala 29:58]
  wire  signProd; // @[MulAddRecFN.scala 98:30]
  wire [13:0] _T_50; // @[MulAddRecFN.scala 101:19]
  wire [13:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  doSubMags; // @[MulAddRecFN.scala 103:30]
  wire [13:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [13:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [12:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _T_57; // @[MulAddRecFN.scala 109:35]
  wire  _T_58; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _T_60; // @[MulAddRecFN.scala 111:60]
  wire  _T_61; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _T_62; // @[MulAddRecFN.scala 115:34]
  wire [7:0] _T_64; // @[MulAddRecFN.scala 115:16]
  wire [7:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [53:0] _T_66; // @[MulAddRecFN.scala 121:16]
  wire [110:0] _T_68; // @[Bitwise.scala 71:12]
  wire [164:0] _T_70; // @[MulAddRecFN.scala 123:11]
  wire [164:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire  _T_74; // @[primitives.scala 121:54]
  wire  _T_76; // @[primitives.scala 121:54]
  wire  _T_78; // @[primitives.scala 121:54]
  wire  _T_80; // @[primitives.scala 121:54]
  wire  _T_82; // @[primitives.scala 121:54]
  wire  _T_84; // @[primitives.scala 121:54]
  wire  _T_86; // @[primitives.scala 121:54]
  wire  _T_88; // @[primitives.scala 121:54]
  wire  _T_90; // @[primitives.scala 121:54]
  wire  _T_92; // @[primitives.scala 121:54]
  wire  _T_94; // @[primitives.scala 121:54]
  wire  _T_96; // @[primitives.scala 121:54]
  wire  _T_98; // @[primitives.scala 121:54]
  wire  _T_100; // @[primitives.scala 124:57]
  wire [6:0] _T_106; // @[primitives.scala 125:20]
  wire [13:0] _T_113; // @[primitives.scala 125:20]
  wire [64:0] _T_115; // @[primitives.scala 77:58]
  wire [7:0] _T_121; // @[Bitwise.scala 102:31]
  wire [7:0] _T_123; // @[Bitwise.scala 102:65]
  wire [7:0] _T_125; // @[Bitwise.scala 102:75]
  wire [7:0] _T_126; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [7:0] _T_131; // @[Bitwise.scala 102:31]
  wire [7:0] _T_133; // @[Bitwise.scala 102:65]
  wire [7:0] _T_135; // @[Bitwise.scala 102:75]
  wire [7:0] _T_136; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 102:31]
  wire [7:0] _T_141; // @[Bitwise.scala 102:31]
  wire [7:0] _T_143; // @[Bitwise.scala 102:65]
  wire [7:0] _T_145; // @[Bitwise.scala 102:75]
  wire [7:0] _T_146; // @[Bitwise.scala 102:39]
  wire [12:0] _T_160; // @[Cat.scala 29:58]
  wire [13:0] _GEN_3; // @[MulAddRecFN.scala 125:68]
  wire [13:0] _T_161; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _T_164; // @[MulAddRecFN.scala 137:39]
  wire  _T_166; // @[MulAddRecFN.scala 137:44]
  wire  _T_168; // @[MulAddRecFN.scala 138:39]
  wire  _T_169; // @[MulAddRecFN.scala 138:44]
  wire  _T_170; // @[MulAddRecFN.scala 136:16]
  wire [161:0] _T_171; // @[Cat.scala 29:58]
  wire [162:0] alignedSigC; // @[Cat.scala 29:58]
  wire  _T_175; // @[common.scala 81:46]
  wire  _T_178; // @[common.scala 81:46]
  wire  _T_179; // @[MulAddRecFN.scala 149:32]
  wire  _T_182; // @[common.scala 81:46]
  wire [13:0] _T_187; // @[MulAddRecFN.scala 161:53]
  wire [13:0] _T_188; // @[MulAddRecFN.scala 161:12]
  assign rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[51:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[51:0]}; // @[Cat.scala 29:58]
  assign rawC_isZero = io_c[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_36 = io_c[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC_isNaN = _T_36 & io_c[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC_sign = io_c[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC_sExp = {1'b0,$signed(io_c[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_sig = {1'h0,~rawC_isZero,io_c[51:0]}; // @[Cat.scala 29:58]
  assign signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_T_50) - 14'sh7c8; // @[MulAddRecFN.scala 101:32]
  assign doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign _GEN_0 = {{1{rawC_sExp[12]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[12:0]; // @[MulAddRecFN.scala 108:42]
  assign _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _T_58 = $signed(sNatCAlignDist) < 14'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50]
  assign _T_60 = posNatCAlignDist <= 13'h35; // @[MulAddRecFN.scala 111:60]
  assign _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 111:23]
  assign _T_62 = posNatCAlignDist < 13'ha1; // @[MulAddRecFN.scala 115:34]
  assign _T_64 = _T_62 ? posNatCAlignDist[7:0] : 8'ha1; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 8'h0 : _T_64; // @[MulAddRecFN.scala 113:12]
  assign _T_66 = doSubMags ? ~rawC_sig : rawC_sig; // @[MulAddRecFN.scala 121:16]
  assign _T_68 = doSubMags ? 111'h7fffffffffffffffffffffffffff : 111'h0; // @[Bitwise.scala 71:12]
  assign _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _T_74 = rawC_sig[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_76 = rawC_sig[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_78 = rawC_sig[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_80 = rawC_sig[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_82 = rawC_sig[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_84 = rawC_sig[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_86 = rawC_sig[27:24] != 4'h0; // @[primitives.scala 121:54]
  assign _T_88 = rawC_sig[31:28] != 4'h0; // @[primitives.scala 121:54]
  assign _T_90 = rawC_sig[35:32] != 4'h0; // @[primitives.scala 121:54]
  assign _T_92 = rawC_sig[39:36] != 4'h0; // @[primitives.scala 121:54]
  assign _T_94 = rawC_sig[43:40] != 4'h0; // @[primitives.scala 121:54]
  assign _T_96 = rawC_sig[47:44] != 4'h0; // @[primitives.scala 121:54]
  assign _T_98 = rawC_sig[51:48] != 4'h0; // @[primitives.scala 121:54]
  assign _T_100 = rawC_sig[53:52] != 2'h0; // @[primitives.scala 124:57]
  assign _T_106 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76,_T_74}; // @[primitives.scala 125:20]
  assign _T_113 = {_T_100,_T_98,_T_96,_T_94,_T_92,_T_90,_T_88,_T_106}; // @[primitives.scala 125:20]
  assign _T_115 = -65'sh10000000000000000 >>> CAlignDist[7:2]; // @[primitives.scala 77:58]
  assign _T_121 = {{4'd0}, _T_115[31:28]}; // @[Bitwise.scala 102:31]
  assign _T_123 = {_T_115[27:24], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_125 = _T_123 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_126 = _T_121 | _T_125; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{2'd0}, _T_126[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_131 = _GEN_1 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_133 = {_T_126[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_135 = _T_133 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_136 = _T_131 | _T_135; // @[Bitwise.scala 102:39]
  assign _GEN_2 = {{1'd0}, _T_136[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_141 = _GEN_2 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_143 = {_T_136[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_145 = _T_143 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_146 = _T_141 | _T_145; // @[Bitwise.scala 102:39]
  assign _T_160 = {_T_146,_T_115[32],_T_115[33],_T_115[34],_T_115[35],_T_115[36]}; // @[Cat.scala 29:58]
  assign _GEN_3 = {{1'd0}, _T_160}; // @[MulAddRecFN.scala 125:68]
  assign _T_161 = _T_113 & _GEN_3; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = _T_161 != 14'h0; // @[MulAddRecFN.scala 133:11]
  assign _T_164 = mainAlignedSigC[2:0] == 3'h7; // @[MulAddRecFN.scala 137:39]
  assign _T_166 = _T_164 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _T_168 = mainAlignedSigC[2:0] != 3'h0; // @[MulAddRecFN.scala 138:39]
  assign _T_169 = _T_168 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign _T_170 = doSubMags ? _T_166 : _T_169; // @[MulAddRecFN.scala 136:16]
  assign _T_171 = mainAlignedSigC[164:3]; // @[Cat.scala 29:58]
  assign alignedSigC = {_T_171,_T_170}; // @[Cat.scala 29:58]
  assign _T_175 = rawA_isNaN & ~rawA_sig[51]; // @[common.scala 81:46]
  assign _T_178 = rawB_isNaN & ~rawB_sig[51]; // @[common.scala 81:46]
  assign _T_179 = _T_175 | _T_178; // @[MulAddRecFN.scala 149:32]
  assign _T_182 = rawC_isNaN & ~rawC_sig[51]; // @[common.scala 81:46]
  assign _T_187 = $signed(sExpAlignedProd) - 14'sh35; // @[MulAddRecFN.scala 161:53]
  assign _T_188 = CIsDominant ? $signed({{1{rawC_sExp[12]}},rawC_sExp}) : $signed(_T_187); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[52:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[52:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[106:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_179 | _T_182; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_4 & ~io_a[61]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[63:61] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_20 & ~io_b[61]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[63:61] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_36 & io_c[61]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_36 & ~io_c[61]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[63:61] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_188[12:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[5:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[161:107]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
endmodule
module MulAddRecFNToRaw_postMul(
  input          io_fromPreMul_isSigNaNAny,
  input          io_fromPreMul_isNaNAOrB,
  input          io_fromPreMul_isInfA,
  input          io_fromPreMul_isZeroA,
  input          io_fromPreMul_isInfB,
  input          io_fromPreMul_isZeroB,
  input          io_fromPreMul_signProd,
  input          io_fromPreMul_isNaNC,
  input          io_fromPreMul_isInfC,
  input          io_fromPreMul_isZeroC,
  input  [12:0]  io_fromPreMul_sExpSum,
  input          io_fromPreMul_doSubMags,
  input          io_fromPreMul_CIsDominant,
  input  [5:0]   io_fromPreMul_CDom_CAlignDist,
  input  [54:0]  io_fromPreMul_highAlignedSigC,
  input          io_fromPreMul_bit0AlignedSigC,
  input  [106:0] io_mulAddResult,
  input  [2:0]   io_roundingMode,
  output         io_invalidExc,
  output         io_rawOut_isNaN,
  output         io_rawOut_isInf,
  output         io_rawOut_isZero,
  output         io_rawOut_sign,
  output [12:0]  io_rawOut_sExp,
  output [55:0]  io_rawOut_sig
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [54:0] _T_2; // @[MulAddRecFN.scala 195:47]
  wire [54:0] _T_3; // @[MulAddRecFN.scala 194:16]
  wire [161:0] sigSum; // @[Cat.scala 29:58]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69]
  wire [12:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [12:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [107:0] _T_14; // @[Cat.scala 29:58]
  wire [107:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _T_17; // @[MulAddRecFN.scala 217:36]
  wire  _T_19; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [170:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [170:0] _T_20; // @[MulAddRecFN.scala 221:24]
  wire [57:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [54:0] _T_22; // @[MulAddRecFN.scala 224:53]
  wire  _T_25; // @[primitives.scala 121:54]
  wire  _T_27; // @[primitives.scala 121:54]
  wire  _T_29; // @[primitives.scala 121:54]
  wire  _T_31; // @[primitives.scala 121:54]
  wire  _T_33; // @[primitives.scala 121:54]
  wire  _T_35; // @[primitives.scala 121:54]
  wire  _T_37; // @[primitives.scala 121:54]
  wire  _T_39; // @[primitives.scala 121:54]
  wire  _T_41; // @[primitives.scala 121:54]
  wire  _T_43; // @[primitives.scala 121:54]
  wire  _T_45; // @[primitives.scala 121:54]
  wire  _T_47; // @[primitives.scala 121:54]
  wire  _T_49; // @[primitives.scala 121:54]
  wire  _T_51; // @[primitives.scala 124:57]
  wire [6:0] _T_57; // @[primitives.scala 125:20]
  wire [13:0] _T_64; // @[primitives.scala 125:20]
  wire [16:0] _T_67; // @[primitives.scala 77:58]
  wire [7:0] _T_73; // @[Bitwise.scala 102:31]
  wire [7:0] _T_75; // @[Bitwise.scala 102:65]
  wire [7:0] _T_77; // @[Bitwise.scala 102:75]
  wire [7:0] _T_78; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 102:31]
  wire [7:0] _T_83; // @[Bitwise.scala 102:31]
  wire [7:0] _T_85; // @[Bitwise.scala 102:65]
  wire [7:0] _T_87; // @[Bitwise.scala 102:75]
  wire [7:0] _T_88; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_3; // @[Bitwise.scala 102:31]
  wire [7:0] _T_93; // @[Bitwise.scala 102:31]
  wire [7:0] _T_95; // @[Bitwise.scala 102:65]
  wire [7:0] _T_97; // @[Bitwise.scala 102:75]
  wire [7:0] _T_98; // @[Bitwise.scala 102:39]
  wire [12:0] _T_112; // @[Cat.scala 29:58]
  wire [13:0] _GEN_4; // @[MulAddRecFN.scala 224:72]
  wire [13:0] _T_113; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire  _T_116; // @[MulAddRecFN.scala 228:32]
  wire  _T_117; // @[MulAddRecFN.scala 228:36]
  wire  _T_118; // @[MulAddRecFN.scala 228:61]
  wire [55:0] CDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [108:0] _GEN_5; // @[MulAddRecFN.scala 238:41]
  wire [108:0] _T_123; // @[MulAddRecFN.scala 238:41]
  wire [108:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  _T_126; // @[primitives.scala 104:54]
  wire  _T_128; // @[primitives.scala 104:54]
  wire  _T_130; // @[primitives.scala 104:54]
  wire  _T_132; // @[primitives.scala 104:54]
  wire  _T_134; // @[primitives.scala 104:54]
  wire  _T_136; // @[primitives.scala 104:54]
  wire  _T_138; // @[primitives.scala 104:54]
  wire  _T_140; // @[primitives.scala 104:54]
  wire  _T_142; // @[primitives.scala 104:54]
  wire  _T_144; // @[primitives.scala 104:54]
  wire  _T_146; // @[primitives.scala 104:54]
  wire  _T_148; // @[primitives.scala 104:54]
  wire  _T_150; // @[primitives.scala 104:54]
  wire  _T_152; // @[primitives.scala 104:54]
  wire  _T_154; // @[primitives.scala 104:54]
  wire  _T_156; // @[primitives.scala 104:54]
  wire  _T_158; // @[primitives.scala 104:54]
  wire  _T_160; // @[primitives.scala 104:54]
  wire  _T_162; // @[primitives.scala 104:54]
  wire  _T_164; // @[primitives.scala 104:54]
  wire  _T_166; // @[primitives.scala 104:54]
  wire  _T_168; // @[primitives.scala 104:54]
  wire  _T_170; // @[primitives.scala 104:54]
  wire  _T_172; // @[primitives.scala 104:54]
  wire  _T_174; // @[primitives.scala 104:54]
  wire  _T_176; // @[primitives.scala 104:54]
  wire  _T_178; // @[primitives.scala 104:54]
  wire  _T_180; // @[primitives.scala 104:54]
  wire  _T_182; // @[primitives.scala 104:54]
  wire  _T_184; // @[primitives.scala 104:54]
  wire  _T_186; // @[primitives.scala 104:54]
  wire  _T_188; // @[primitives.scala 104:54]
  wire  _T_190; // @[primitives.scala 104:54]
  wire  _T_192; // @[primitives.scala 104:54]
  wire  _T_194; // @[primitives.scala 104:54]
  wire  _T_196; // @[primitives.scala 104:54]
  wire  _T_198; // @[primitives.scala 104:54]
  wire  _T_200; // @[primitives.scala 104:54]
  wire  _T_202; // @[primitives.scala 104:54]
  wire  _T_204; // @[primitives.scala 104:54]
  wire  _T_206; // @[primitives.scala 104:54]
  wire  _T_208; // @[primitives.scala 104:54]
  wire  _T_210; // @[primitives.scala 104:54]
  wire  _T_212; // @[primitives.scala 104:54]
  wire  _T_214; // @[primitives.scala 104:54]
  wire  _T_216; // @[primitives.scala 104:54]
  wire  _T_218; // @[primitives.scala 104:54]
  wire  _T_220; // @[primitives.scala 104:54]
  wire  _T_222; // @[primitives.scala 104:54]
  wire  _T_224; // @[primitives.scala 104:54]
  wire  _T_226; // @[primitives.scala 104:54]
  wire  _T_228; // @[primitives.scala 104:54]
  wire  _T_230; // @[primitives.scala 104:54]
  wire  _T_232; // @[primitives.scala 104:54]
  wire [5:0] _T_239; // @[primitives.scala 108:20]
  wire [12:0] _T_246; // @[primitives.scala 108:20]
  wire [6:0] _T_252; // @[primitives.scala 108:20]
  wire [26:0] _T_260; // @[primitives.scala 108:20]
  wire [6:0] _T_266; // @[primitives.scala 108:20]
  wire [13:0] _T_273; // @[primitives.scala 108:20]
  wire [6:0] _T_279; // @[primitives.scala 108:20]
  wire [54:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [5:0] _T_343; // @[Mux.scala 47:69]
  wire [5:0] _T_344; // @[Mux.scala 47:69]
  wire [5:0] _T_345; // @[Mux.scala 47:69]
  wire [5:0] _T_346; // @[Mux.scala 47:69]
  wire [5:0] _T_347; // @[Mux.scala 47:69]
  wire [5:0] _T_348; // @[Mux.scala 47:69]
  wire [5:0] _T_349; // @[Mux.scala 47:69]
  wire [5:0] _T_350; // @[Mux.scala 47:69]
  wire [5:0] _T_351; // @[Mux.scala 47:69]
  wire [5:0] _T_352; // @[Mux.scala 47:69]
  wire [5:0] _T_353; // @[Mux.scala 47:69]
  wire [5:0] _T_354; // @[Mux.scala 47:69]
  wire [5:0] _T_355; // @[Mux.scala 47:69]
  wire [5:0] _T_356; // @[Mux.scala 47:69]
  wire [5:0] _T_357; // @[Mux.scala 47:69]
  wire [5:0] _T_358; // @[Mux.scala 47:69]
  wire [5:0] _T_359; // @[Mux.scala 47:69]
  wire [5:0] _T_360; // @[Mux.scala 47:69]
  wire [5:0] _T_361; // @[Mux.scala 47:69]
  wire [5:0] _T_362; // @[Mux.scala 47:69]
  wire [5:0] _T_363; // @[Mux.scala 47:69]
  wire [5:0] _T_364; // @[Mux.scala 47:69]
  wire [5:0] _T_365; // @[Mux.scala 47:69]
  wire [5:0] _T_366; // @[Mux.scala 47:69]
  wire [5:0] _T_367; // @[Mux.scala 47:69]
  wire [5:0] _T_368; // @[Mux.scala 47:69]
  wire [5:0] _T_369; // @[Mux.scala 47:69]
  wire [5:0] _T_370; // @[Mux.scala 47:69]
  wire [5:0] _T_371; // @[Mux.scala 47:69]
  wire [5:0] _T_372; // @[Mux.scala 47:69]
  wire [5:0] _T_373; // @[Mux.scala 47:69]
  wire [5:0] _T_374; // @[Mux.scala 47:69]
  wire [5:0] _T_375; // @[Mux.scala 47:69]
  wire [5:0] _T_376; // @[Mux.scala 47:69]
  wire [5:0] _T_377; // @[Mux.scala 47:69]
  wire [5:0] _T_378; // @[Mux.scala 47:69]
  wire [5:0] _T_379; // @[Mux.scala 47:69]
  wire [5:0] _T_380; // @[Mux.scala 47:69]
  wire [5:0] _T_381; // @[Mux.scala 47:69]
  wire [5:0] _T_382; // @[Mux.scala 47:69]
  wire [5:0] _T_383; // @[Mux.scala 47:69]
  wire [5:0] _T_384; // @[Mux.scala 47:69]
  wire [5:0] _T_385; // @[Mux.scala 47:69]
  wire [5:0] _T_386; // @[Mux.scala 47:69]
  wire [5:0] _T_387; // @[Mux.scala 47:69]
  wire [5:0] _T_388; // @[Mux.scala 47:69]
  wire [5:0] _T_389; // @[Mux.scala 47:69]
  wire [5:0] _T_390; // @[Mux.scala 47:69]
  wire [5:0] _T_391; // @[Mux.scala 47:69]
  wire [5:0] _T_392; // @[Mux.scala 47:69]
  wire [5:0] _T_393; // @[Mux.scala 47:69]
  wire [5:0] _T_394; // @[Mux.scala 47:69]
  wire [5:0] _T_395; // @[Mux.scala 47:69]
  wire [5:0] notCDom_normDistReduced2; // @[Mux.scala 47:69]
  wire [6:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [7:0] _T_396; // @[MulAddRecFN.scala 243:69]
  wire [12:0] _GEN_6; // @[MulAddRecFN.scala 243:46]
  wire [12:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [235:0] _GEN_7; // @[MulAddRecFN.scala 245:27]
  wire [235:0] _T_399; // @[MulAddRecFN.scala 245:27]
  wire [57:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  _T_404; // @[primitives.scala 104:54]
  wire  _T_406; // @[primitives.scala 104:54]
  wire  _T_408; // @[primitives.scala 104:54]
  wire  _T_410; // @[primitives.scala 104:54]
  wire  _T_412; // @[primitives.scala 104:54]
  wire  _T_414; // @[primitives.scala 104:54]
  wire  _T_416; // @[primitives.scala 104:54]
  wire  _T_418; // @[primitives.scala 104:54]
  wire  _T_420; // @[primitives.scala 104:54]
  wire  _T_422; // @[primitives.scala 104:54]
  wire  _T_424; // @[primitives.scala 104:54]
  wire  _T_426; // @[primitives.scala 104:54]
  wire  _T_428; // @[primitives.scala 104:54]
  wire [6:0] _T_436; // @[primitives.scala 108:20]
  wire [13:0] _T_443; // @[primitives.scala 108:20]
  wire [32:0] _T_446; // @[primitives.scala 77:58]
  wire [7:0] _T_452; // @[Bitwise.scala 102:31]
  wire [7:0] _T_454; // @[Bitwise.scala 102:65]
  wire [7:0] _T_456; // @[Bitwise.scala 102:75]
  wire [7:0] _T_457; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_8; // @[Bitwise.scala 102:31]
  wire [7:0] _T_462; // @[Bitwise.scala 102:31]
  wire [7:0] _T_464; // @[Bitwise.scala 102:65]
  wire [7:0] _T_466; // @[Bitwise.scala 102:75]
  wire [7:0] _T_467; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_9; // @[Bitwise.scala 102:31]
  wire [7:0] _T_472; // @[Bitwise.scala 102:31]
  wire [7:0] _T_474; // @[Bitwise.scala 102:65]
  wire [7:0] _T_476; // @[Bitwise.scala 102:75]
  wire [7:0] _T_477; // @[Bitwise.scala 102:39]
  wire [12:0] _T_491; // @[Cat.scala 29:58]
  wire [13:0] _GEN_10; // @[MulAddRecFN.scala 249:78]
  wire [13:0] _T_492; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire  _T_495; // @[MulAddRecFN.scala 254:35]
  wire  _T_496; // @[MulAddRecFN.scala 254:39]
  wire [55:0] notCDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _T_498; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _T_499; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _T_500; // @[MulAddRecFN.scala 274:31]
  wire  _T_501; // @[MulAddRecFN.scala 273:35]
  wire  _T_502; // @[MulAddRecFN.scala 275:32]
  wire  _T_503; // @[MulAddRecFN.scala 274:57]
  wire  _T_506; // @[MulAddRecFN.scala 276:36]
  wire  _T_507; // @[MulAddRecFN.scala 277:61]
  wire  _T_508; // @[MulAddRecFN.scala 278:35]
  wire  _T_512; // @[MulAddRecFN.scala 285:42]
  wire  _T_514; // @[MulAddRecFN.scala 287:27]
  wire  _T_515; // @[MulAddRecFN.scala 288:31]
  wire  _T_516; // @[MulAddRecFN.scala 287:54]
  wire  _T_518; // @[MulAddRecFN.scala 289:26]
  wire  _T_519; // @[MulAddRecFN.scala 289:48]
  wire  _T_520; // @[MulAddRecFN.scala 290:36]
  wire  _T_521; // @[MulAddRecFN.scala 288:43]
  wire  _T_522; // @[MulAddRecFN.scala 291:26]
  wire  _T_523; // @[MulAddRecFN.scala 292:37]
  wire  _T_524; // @[MulAddRecFN.scala 291:46]
  wire  _T_525; // @[MulAddRecFN.scala 290:48]
  wire  _T_528; // @[MulAddRecFN.scala 293:28]
  wire  _T_529; // @[MulAddRecFN.scala 294:17]
  wire  _T_530; // @[MulAddRecFN.scala 293:49]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 55'h1; // @[MulAddRecFN.scala 195:47]
  assign _T_3 = io_mulAddResult[106] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum = {_T_3,io_mulAddResult[105:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{11{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[54:53],sigSum[159:55]}; // @[Cat.scala 29:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[161:54] : _T_14; // @[MulAddRecFN.scala 207:12]
  assign _T_17 = ~sigSum[53:1] != 53'h0; // @[MulAddRecFN.scala 217:36]
  assign _T_19 = sigSum[54:1] != 54'h0; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{63'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _T_20[107:50]; // @[MulAddRecFN.scala 221:56]
  assign _T_22 = {CDom_absSigSum[52:0], 2'h0}; // @[MulAddRecFN.scala 224:53]
  assign _T_25 = _T_22[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_27 = _T_22[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_29 = _T_22[11:8] != 4'h0; // @[primitives.scala 121:54]
  assign _T_31 = _T_22[15:12] != 4'h0; // @[primitives.scala 121:54]
  assign _T_33 = _T_22[19:16] != 4'h0; // @[primitives.scala 121:54]
  assign _T_35 = _T_22[23:20] != 4'h0; // @[primitives.scala 121:54]
  assign _T_37 = _T_22[27:24] != 4'h0; // @[primitives.scala 121:54]
  assign _T_39 = _T_22[31:28] != 4'h0; // @[primitives.scala 121:54]
  assign _T_41 = _T_22[35:32] != 4'h0; // @[primitives.scala 121:54]
  assign _T_43 = _T_22[39:36] != 4'h0; // @[primitives.scala 121:54]
  assign _T_45 = _T_22[43:40] != 4'h0; // @[primitives.scala 121:54]
  assign _T_47 = _T_22[47:44] != 4'h0; // @[primitives.scala 121:54]
  assign _T_49 = _T_22[51:48] != 4'h0; // @[primitives.scala 121:54]
  assign _T_51 = _T_22[54:52] != 3'h0; // @[primitives.scala 124:57]
  assign _T_57 = {_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25}; // @[primitives.scala 125:20]
  assign _T_64 = {_T_51,_T_49,_T_47,_T_45,_T_43,_T_41,_T_39,_T_57}; // @[primitives.scala 125:20]
  assign _T_67 = -17'sh10000 >>> ~io_fromPreMul_CDom_CAlignDist[5:2]; // @[primitives.scala 77:58]
  assign _T_73 = {{4'd0}, _T_67[8:5]}; // @[Bitwise.scala 102:31]
  assign _T_75 = {_T_67[4:1], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_77 = _T_75 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_78 = _T_73 | _T_77; // @[Bitwise.scala 102:39]
  assign _GEN_2 = {{2'd0}, _T_78[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_83 = _GEN_2 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_85 = {_T_78[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_87 = _T_85 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_88 = _T_83 | _T_87; // @[Bitwise.scala 102:39]
  assign _GEN_3 = {{1'd0}, _T_88[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_93 = _GEN_3 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_95 = {_T_88[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_97 = _T_95 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_98 = _T_93 | _T_97; // @[Bitwise.scala 102:39]
  assign _T_112 = {_T_98,_T_67[9],_T_67[10],_T_67[11],_T_67[12],_T_67[13]}; // @[Cat.scala 29:58]
  assign _GEN_4 = {{1'd0}, _T_112}; // @[MulAddRecFN.scala 224:72]
  assign _T_113 = _T_64 & _GEN_4; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = _T_113 != 14'h0; // @[MulAddRecFN.scala 225:73]
  assign _T_116 = CDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 228:32]
  assign _T_117 = _T_116 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign _T_118 = _T_117 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_mainSig[57:3],_T_118}; // @[Cat.scala 29:58]
  assign notCDom_signSigSum = sigSum[109]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_5 = {{108'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _T_123 = sigSum[108:0] + _GEN_5; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[108:0] : _T_123; // @[MulAddRecFN.scala 236:12]
  assign _T_126 = notCDom_absSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_128 = notCDom_absSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_130 = notCDom_absSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_132 = notCDom_absSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_134 = notCDom_absSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_136 = notCDom_absSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_138 = notCDom_absSigSum[13:12] != 2'h0; // @[primitives.scala 104:54]
  assign _T_140 = notCDom_absSigSum[15:14] != 2'h0; // @[primitives.scala 104:54]
  assign _T_142 = notCDom_absSigSum[17:16] != 2'h0; // @[primitives.scala 104:54]
  assign _T_144 = notCDom_absSigSum[19:18] != 2'h0; // @[primitives.scala 104:54]
  assign _T_146 = notCDom_absSigSum[21:20] != 2'h0; // @[primitives.scala 104:54]
  assign _T_148 = notCDom_absSigSum[23:22] != 2'h0; // @[primitives.scala 104:54]
  assign _T_150 = notCDom_absSigSum[25:24] != 2'h0; // @[primitives.scala 104:54]
  assign _T_152 = notCDom_absSigSum[27:26] != 2'h0; // @[primitives.scala 104:54]
  assign _T_154 = notCDom_absSigSum[29:28] != 2'h0; // @[primitives.scala 104:54]
  assign _T_156 = notCDom_absSigSum[31:30] != 2'h0; // @[primitives.scala 104:54]
  assign _T_158 = notCDom_absSigSum[33:32] != 2'h0; // @[primitives.scala 104:54]
  assign _T_160 = notCDom_absSigSum[35:34] != 2'h0; // @[primitives.scala 104:54]
  assign _T_162 = notCDom_absSigSum[37:36] != 2'h0; // @[primitives.scala 104:54]
  assign _T_164 = notCDom_absSigSum[39:38] != 2'h0; // @[primitives.scala 104:54]
  assign _T_166 = notCDom_absSigSum[41:40] != 2'h0; // @[primitives.scala 104:54]
  assign _T_168 = notCDom_absSigSum[43:42] != 2'h0; // @[primitives.scala 104:54]
  assign _T_170 = notCDom_absSigSum[45:44] != 2'h0; // @[primitives.scala 104:54]
  assign _T_172 = notCDom_absSigSum[47:46] != 2'h0; // @[primitives.scala 104:54]
  assign _T_174 = notCDom_absSigSum[49:48] != 2'h0; // @[primitives.scala 104:54]
  assign _T_176 = notCDom_absSigSum[51:50] != 2'h0; // @[primitives.scala 104:54]
  assign _T_178 = notCDom_absSigSum[53:52] != 2'h0; // @[primitives.scala 104:54]
  assign _T_180 = notCDom_absSigSum[55:54] != 2'h0; // @[primitives.scala 104:54]
  assign _T_182 = notCDom_absSigSum[57:56] != 2'h0; // @[primitives.scala 104:54]
  assign _T_184 = notCDom_absSigSum[59:58] != 2'h0; // @[primitives.scala 104:54]
  assign _T_186 = notCDom_absSigSum[61:60] != 2'h0; // @[primitives.scala 104:54]
  assign _T_188 = notCDom_absSigSum[63:62] != 2'h0; // @[primitives.scala 104:54]
  assign _T_190 = notCDom_absSigSum[65:64] != 2'h0; // @[primitives.scala 104:54]
  assign _T_192 = notCDom_absSigSum[67:66] != 2'h0; // @[primitives.scala 104:54]
  assign _T_194 = notCDom_absSigSum[69:68] != 2'h0; // @[primitives.scala 104:54]
  assign _T_196 = notCDom_absSigSum[71:70] != 2'h0; // @[primitives.scala 104:54]
  assign _T_198 = notCDom_absSigSum[73:72] != 2'h0; // @[primitives.scala 104:54]
  assign _T_200 = notCDom_absSigSum[75:74] != 2'h0; // @[primitives.scala 104:54]
  assign _T_202 = notCDom_absSigSum[77:76] != 2'h0; // @[primitives.scala 104:54]
  assign _T_204 = notCDom_absSigSum[79:78] != 2'h0; // @[primitives.scala 104:54]
  assign _T_206 = notCDom_absSigSum[81:80] != 2'h0; // @[primitives.scala 104:54]
  assign _T_208 = notCDom_absSigSum[83:82] != 2'h0; // @[primitives.scala 104:54]
  assign _T_210 = notCDom_absSigSum[85:84] != 2'h0; // @[primitives.scala 104:54]
  assign _T_212 = notCDom_absSigSum[87:86] != 2'h0; // @[primitives.scala 104:54]
  assign _T_214 = notCDom_absSigSum[89:88] != 2'h0; // @[primitives.scala 104:54]
  assign _T_216 = notCDom_absSigSum[91:90] != 2'h0; // @[primitives.scala 104:54]
  assign _T_218 = notCDom_absSigSum[93:92] != 2'h0; // @[primitives.scala 104:54]
  assign _T_220 = notCDom_absSigSum[95:94] != 2'h0; // @[primitives.scala 104:54]
  assign _T_222 = notCDom_absSigSum[97:96] != 2'h0; // @[primitives.scala 104:54]
  assign _T_224 = notCDom_absSigSum[99:98] != 2'h0; // @[primitives.scala 104:54]
  assign _T_226 = notCDom_absSigSum[101:100] != 2'h0; // @[primitives.scala 104:54]
  assign _T_228 = notCDom_absSigSum[103:102] != 2'h0; // @[primitives.scala 104:54]
  assign _T_230 = notCDom_absSigSum[105:104] != 2'h0; // @[primitives.scala 104:54]
  assign _T_232 = notCDom_absSigSum[107:106] != 2'h0; // @[primitives.scala 104:54]
  assign _T_239 = {_T_136,_T_134,_T_132,_T_130,_T_128,_T_126}; // @[primitives.scala 108:20]
  assign _T_246 = {_T_150,_T_148,_T_146,_T_144,_T_142,_T_140,_T_138,_T_239}; // @[primitives.scala 108:20]
  assign _T_252 = {_T_164,_T_162,_T_160,_T_158,_T_156,_T_154,_T_152}; // @[primitives.scala 108:20]
  assign _T_260 = {_T_178,_T_176,_T_174,_T_172,_T_170,_T_168,_T_166,_T_252,_T_246}; // @[primitives.scala 108:20]
  assign _T_266 = {_T_192,_T_190,_T_188,_T_186,_T_184,_T_182,_T_180}; // @[primitives.scala 108:20]
  assign _T_273 = {_T_206,_T_204,_T_202,_T_200,_T_198,_T_196,_T_194,_T_266}; // @[primitives.scala 108:20]
  assign _T_279 = {_T_220,_T_218,_T_216,_T_214,_T_212,_T_210,_T_208}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {notCDom_absSigSum[108],_T_232,_T_230,_T_228,_T_226,_T_224,_T_222,_T_279,_T_273,_T_260}; // @[primitives.scala 108:20]
  assign _T_343 = notCDom_reduced2AbsSigSum[1] ? 6'h35 : 6'h36; // @[Mux.scala 47:69]
  assign _T_344 = notCDom_reduced2AbsSigSum[2] ? 6'h34 : _T_343; // @[Mux.scala 47:69]
  assign _T_345 = notCDom_reduced2AbsSigSum[3] ? 6'h33 : _T_344; // @[Mux.scala 47:69]
  assign _T_346 = notCDom_reduced2AbsSigSum[4] ? 6'h32 : _T_345; // @[Mux.scala 47:69]
  assign _T_347 = notCDom_reduced2AbsSigSum[5] ? 6'h31 : _T_346; // @[Mux.scala 47:69]
  assign _T_348 = notCDom_reduced2AbsSigSum[6] ? 6'h30 : _T_347; // @[Mux.scala 47:69]
  assign _T_349 = notCDom_reduced2AbsSigSum[7] ? 6'h2f : _T_348; // @[Mux.scala 47:69]
  assign _T_350 = notCDom_reduced2AbsSigSum[8] ? 6'h2e : _T_349; // @[Mux.scala 47:69]
  assign _T_351 = notCDom_reduced2AbsSigSum[9] ? 6'h2d : _T_350; // @[Mux.scala 47:69]
  assign _T_352 = notCDom_reduced2AbsSigSum[10] ? 6'h2c : _T_351; // @[Mux.scala 47:69]
  assign _T_353 = notCDom_reduced2AbsSigSum[11] ? 6'h2b : _T_352; // @[Mux.scala 47:69]
  assign _T_354 = notCDom_reduced2AbsSigSum[12] ? 6'h2a : _T_353; // @[Mux.scala 47:69]
  assign _T_355 = notCDom_reduced2AbsSigSum[13] ? 6'h29 : _T_354; // @[Mux.scala 47:69]
  assign _T_356 = notCDom_reduced2AbsSigSum[14] ? 6'h28 : _T_355; // @[Mux.scala 47:69]
  assign _T_357 = notCDom_reduced2AbsSigSum[15] ? 6'h27 : _T_356; // @[Mux.scala 47:69]
  assign _T_358 = notCDom_reduced2AbsSigSum[16] ? 6'h26 : _T_357; // @[Mux.scala 47:69]
  assign _T_359 = notCDom_reduced2AbsSigSum[17] ? 6'h25 : _T_358; // @[Mux.scala 47:69]
  assign _T_360 = notCDom_reduced2AbsSigSum[18] ? 6'h24 : _T_359; // @[Mux.scala 47:69]
  assign _T_361 = notCDom_reduced2AbsSigSum[19] ? 6'h23 : _T_360; // @[Mux.scala 47:69]
  assign _T_362 = notCDom_reduced2AbsSigSum[20] ? 6'h22 : _T_361; // @[Mux.scala 47:69]
  assign _T_363 = notCDom_reduced2AbsSigSum[21] ? 6'h21 : _T_362; // @[Mux.scala 47:69]
  assign _T_364 = notCDom_reduced2AbsSigSum[22] ? 6'h20 : _T_363; // @[Mux.scala 47:69]
  assign _T_365 = notCDom_reduced2AbsSigSum[23] ? 6'h1f : _T_364; // @[Mux.scala 47:69]
  assign _T_366 = notCDom_reduced2AbsSigSum[24] ? 6'h1e : _T_365; // @[Mux.scala 47:69]
  assign _T_367 = notCDom_reduced2AbsSigSum[25] ? 6'h1d : _T_366; // @[Mux.scala 47:69]
  assign _T_368 = notCDom_reduced2AbsSigSum[26] ? 6'h1c : _T_367; // @[Mux.scala 47:69]
  assign _T_369 = notCDom_reduced2AbsSigSum[27] ? 6'h1b : _T_368; // @[Mux.scala 47:69]
  assign _T_370 = notCDom_reduced2AbsSigSum[28] ? 6'h1a : _T_369; // @[Mux.scala 47:69]
  assign _T_371 = notCDom_reduced2AbsSigSum[29] ? 6'h19 : _T_370; // @[Mux.scala 47:69]
  assign _T_372 = notCDom_reduced2AbsSigSum[30] ? 6'h18 : _T_371; // @[Mux.scala 47:69]
  assign _T_373 = notCDom_reduced2AbsSigSum[31] ? 6'h17 : _T_372; // @[Mux.scala 47:69]
  assign _T_374 = notCDom_reduced2AbsSigSum[32] ? 6'h16 : _T_373; // @[Mux.scala 47:69]
  assign _T_375 = notCDom_reduced2AbsSigSum[33] ? 6'h15 : _T_374; // @[Mux.scala 47:69]
  assign _T_376 = notCDom_reduced2AbsSigSum[34] ? 6'h14 : _T_375; // @[Mux.scala 47:69]
  assign _T_377 = notCDom_reduced2AbsSigSum[35] ? 6'h13 : _T_376; // @[Mux.scala 47:69]
  assign _T_378 = notCDom_reduced2AbsSigSum[36] ? 6'h12 : _T_377; // @[Mux.scala 47:69]
  assign _T_379 = notCDom_reduced2AbsSigSum[37] ? 6'h11 : _T_378; // @[Mux.scala 47:69]
  assign _T_380 = notCDom_reduced2AbsSigSum[38] ? 6'h10 : _T_379; // @[Mux.scala 47:69]
  assign _T_381 = notCDom_reduced2AbsSigSum[39] ? 6'hf : _T_380; // @[Mux.scala 47:69]
  assign _T_382 = notCDom_reduced2AbsSigSum[40] ? 6'he : _T_381; // @[Mux.scala 47:69]
  assign _T_383 = notCDom_reduced2AbsSigSum[41] ? 6'hd : _T_382; // @[Mux.scala 47:69]
  assign _T_384 = notCDom_reduced2AbsSigSum[42] ? 6'hc : _T_383; // @[Mux.scala 47:69]
  assign _T_385 = notCDom_reduced2AbsSigSum[43] ? 6'hb : _T_384; // @[Mux.scala 47:69]
  assign _T_386 = notCDom_reduced2AbsSigSum[44] ? 6'ha : _T_385; // @[Mux.scala 47:69]
  assign _T_387 = notCDom_reduced2AbsSigSum[45] ? 6'h9 : _T_386; // @[Mux.scala 47:69]
  assign _T_388 = notCDom_reduced2AbsSigSum[46] ? 6'h8 : _T_387; // @[Mux.scala 47:69]
  assign _T_389 = notCDom_reduced2AbsSigSum[47] ? 6'h7 : _T_388; // @[Mux.scala 47:69]
  assign _T_390 = notCDom_reduced2AbsSigSum[48] ? 6'h6 : _T_389; // @[Mux.scala 47:69]
  assign _T_391 = notCDom_reduced2AbsSigSum[49] ? 6'h5 : _T_390; // @[Mux.scala 47:69]
  assign _T_392 = notCDom_reduced2AbsSigSum[50] ? 6'h4 : _T_391; // @[Mux.scala 47:69]
  assign _T_393 = notCDom_reduced2AbsSigSum[51] ? 6'h3 : _T_392; // @[Mux.scala 47:69]
  assign _T_394 = notCDom_reduced2AbsSigSum[52] ? 6'h2 : _T_393; // @[Mux.scala 47:69]
  assign _T_395 = notCDom_reduced2AbsSigSum[53] ? 6'h1 : _T_394; // @[Mux.scala 47:69]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[54] ? 6'h0 : _T_395; // @[Mux.scala 47:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _T_396 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_6 = {{5{_T_396[7]}},_T_396}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_6); // @[MulAddRecFN.scala 243:46]
  assign _GEN_7 = {{127'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _T_399 = _GEN_7 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _T_399[109:52]; // @[MulAddRecFN.scala 245:50]
  assign _T_404 = notCDom_reduced2AbsSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_406 = notCDom_reduced2AbsSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_408 = notCDom_reduced2AbsSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_410 = notCDom_reduced2AbsSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_412 = notCDom_reduced2AbsSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_414 = notCDom_reduced2AbsSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_416 = notCDom_reduced2AbsSigSum[13:12] != 2'h0; // @[primitives.scala 104:54]
  assign _T_418 = notCDom_reduced2AbsSigSum[15:14] != 2'h0; // @[primitives.scala 104:54]
  assign _T_420 = notCDom_reduced2AbsSigSum[17:16] != 2'h0; // @[primitives.scala 104:54]
  assign _T_422 = notCDom_reduced2AbsSigSum[19:18] != 2'h0; // @[primitives.scala 104:54]
  assign _T_424 = notCDom_reduced2AbsSigSum[21:20] != 2'h0; // @[primitives.scala 104:54]
  assign _T_426 = notCDom_reduced2AbsSigSum[23:22] != 2'h0; // @[primitives.scala 104:54]
  assign _T_428 = notCDom_reduced2AbsSigSum[25:24] != 2'h0; // @[primitives.scala 104:54]
  assign _T_436 = {_T_416,_T_414,_T_412,_T_410,_T_408,_T_406,_T_404}; // @[primitives.scala 108:20]
  assign _T_443 = {notCDom_reduced2AbsSigSum[26],_T_428,_T_426,_T_424,_T_422,_T_420,_T_418,_T_436}; // @[primitives.scala 108:20]
  assign _T_446 = -33'sh100000000 >>> ~notCDom_normDistReduced2[5:1]; // @[primitives.scala 77:58]
  assign _T_452 = {{4'd0}, _T_446[8:5]}; // @[Bitwise.scala 102:31]
  assign _T_454 = {_T_446[4:1], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_456 = _T_454 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_457 = _T_452 | _T_456; // @[Bitwise.scala 102:39]
  assign _GEN_8 = {{2'd0}, _T_457[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_462 = _GEN_8 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_464 = {_T_457[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_466 = _T_464 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_467 = _T_462 | _T_466; // @[Bitwise.scala 102:39]
  assign _GEN_9 = {{1'd0}, _T_467[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_472 = _GEN_9 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_474 = {_T_467[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_476 = _T_474 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_477 = _T_472 | _T_476; // @[Bitwise.scala 102:39]
  assign _T_491 = {_T_477,_T_446[9],_T_446[10],_T_446[11],_T_446[12],_T_446[13]}; // @[Cat.scala 29:58]
  assign _GEN_10 = {{1'd0}, _T_491}; // @[MulAddRecFN.scala 249:78]
  assign _T_492 = _T_443 & _GEN_10; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = _T_492 != 14'h0; // @[MulAddRecFN.scala 251:11]
  assign _T_495 = notCDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 254:35]
  assign _T_496 = _T_495 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_mainSig[57:3],_T_496}; // @[Cat.scala 29:58]
  assign notCDom_completeCancellation = notCDom_sig[55:54] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _T_498 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_498; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _T_499 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _T_499 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _T_500 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _T_501 = io_fromPreMul_isSigNaNAny | _T_500; // @[MulAddRecFN.scala 273:35]
  assign _T_502 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _T_503 = _T_501 | _T_502; // @[MulAddRecFN.scala 274:57]
  assign _T_506 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _T_507 = _T_506 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _T_508 = _T_507 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _T_512 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _T_514 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _T_515 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _T_516 = _T_514 | _T_515; // @[MulAddRecFN.scala 287:54]
  assign _T_518 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _T_519 = _T_518 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _T_520 = _T_519 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _T_521 = _T_516 | _T_520; // @[MulAddRecFN.scala 288:43]
  assign _T_522 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _T_523 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _T_524 = _T_522 & _T_523; // @[MulAddRecFN.scala 291:46]
  assign _T_525 = _T_521 | _T_524; // @[MulAddRecFN.scala 290:48]
  assign _T_528 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _T_529 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _T_530 = _T_528 & _T_529; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_503 | _T_508; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_512; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_525 | _T_530; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  _T_5; // @[primitives.scala 57:25]
  wire  _T_7; // @[primitives.scala 57:25]
  wire  _T_9; // @[primitives.scala 57:25]
  wire  _T_11; // @[primitives.scala 57:25]
  wire  _T_13; // @[primitives.scala 57:25]
  wire  _T_15; // @[primitives.scala 57:25]
  wire [5:0] _T_16; // @[primitives.scala 58:26]
  wire [64:0] _T_17; // @[primitives.scala 77:58]
  wire [31:0] _T_23; // @[Bitwise.scala 102:31]
  wire [31:0] _T_25; // @[Bitwise.scala 102:65]
  wire [31:0] _T_27; // @[Bitwise.scala 102:75]
  wire [31:0] _T_28; // @[Bitwise.scala 102:39]
  wire [31:0] _GEN_0; // @[Bitwise.scala 102:31]
  wire [31:0] _T_33; // @[Bitwise.scala 102:31]
  wire [31:0] _T_35; // @[Bitwise.scala 102:65]
  wire [31:0] _T_37; // @[Bitwise.scala 102:75]
  wire [31:0] _T_38; // @[Bitwise.scala 102:39]
  wire [31:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [31:0] _T_43; // @[Bitwise.scala 102:31]
  wire [31:0] _T_45; // @[Bitwise.scala 102:65]
  wire [31:0] _T_47; // @[Bitwise.scala 102:75]
  wire [31:0] _T_48; // @[Bitwise.scala 102:39]
  wire [31:0] _GEN_2; // @[Bitwise.scala 102:31]
  wire [31:0] _T_53; // @[Bitwise.scala 102:31]
  wire [31:0] _T_55; // @[Bitwise.scala 102:65]
  wire [31:0] _T_57; // @[Bitwise.scala 102:75]
  wire [31:0] _T_58; // @[Bitwise.scala 102:39]
  wire [31:0] _GEN_3; // @[Bitwise.scala 102:31]
  wire [31:0] _T_63; // @[Bitwise.scala 102:31]
  wire [31:0] _T_65; // @[Bitwise.scala 102:65]
  wire [31:0] _T_67; // @[Bitwise.scala 102:75]
  wire [31:0] _T_68; // @[Bitwise.scala 102:39]
  wire [15:0] _T_74; // @[Bitwise.scala 102:31]
  wire [15:0] _T_76; // @[Bitwise.scala 102:65]
  wire [15:0] _T_78; // @[Bitwise.scala 102:75]
  wire [15:0] _T_79; // @[Bitwise.scala 102:39]
  wire [15:0] _GEN_4; // @[Bitwise.scala 102:31]
  wire [15:0] _T_84; // @[Bitwise.scala 102:31]
  wire [15:0] _T_86; // @[Bitwise.scala 102:65]
  wire [15:0] _T_88; // @[Bitwise.scala 102:75]
  wire [15:0] _T_89; // @[Bitwise.scala 102:39]
  wire [15:0] _GEN_5; // @[Bitwise.scala 102:31]
  wire [15:0] _T_94; // @[Bitwise.scala 102:31]
  wire [15:0] _T_96; // @[Bitwise.scala 102:65]
  wire [15:0] _T_98; // @[Bitwise.scala 102:75]
  wire [15:0] _T_99; // @[Bitwise.scala 102:39]
  wire [15:0] _GEN_6; // @[Bitwise.scala 102:31]
  wire [15:0] _T_104; // @[Bitwise.scala 102:31]
  wire [15:0] _T_106; // @[Bitwise.scala 102:65]
  wire [15:0] _T_108; // @[Bitwise.scala 102:75]
  wire [15:0] _T_109; // @[Bitwise.scala 102:39]
  wire [50:0] _T_118; // @[Cat.scala 29:58]
  wire [50:0] _T_120; // @[primitives.scala 74:21]
  wire [50:0] _T_123; // @[primitives.scala 74:21]
  wire [50:0] _T_126; // @[primitives.scala 74:21]
  wire [50:0] _T_129; // @[primitives.scala 74:21]
  wire [53:0] _T_131; // @[Cat.scala 29:58]
  wire [2:0] _T_147; // @[Cat.scala 29:58]
  wire [2:0] _T_148; // @[primitives.scala 61:24]
  wire [2:0] _T_149; // @[primitives.scala 61:24]
  wire [2:0] _T_150; // @[primitives.scala 61:24]
  wire [2:0] _T_151; // @[primitives.scala 61:24]
  wire [53:0] _T_152; // @[primitives.scala 66:24]
  wire [53:0] _T_153; // @[primitives.scala 61:24]
  wire [53:0] _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [53:0] _T_154; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [55:0] _T_155; // @[Cat.scala 29:58]
  wire [55:0] _T_157; // @[Cat.scala 29:58]
  wire [55:0] _T_159; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [55:0] _T_160; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _T_162; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_163; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_164; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_165; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_166; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_167; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_168; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _T_169; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _T_171; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [54:0] _T_176; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _T_178; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _T_180; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_182; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [54:0] _T_184; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_8; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_185; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_9; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] _T_189; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_194; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_199; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _T_201; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _T_203; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_204; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _T_206; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_207; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_208; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  _T_211; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _T_212; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_213; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_214; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_217; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _T_218; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_222; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _T_224; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_225; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_226; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_227; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_229; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _T_234; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_236; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_238; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_239; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_241; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_242; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [11:0] _T_243; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _T_245; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [11:0] _T_247; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [11:0] _T_249; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [11:0] _T_250; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [11:0] _T_252; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [11:0] _T_253; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [11:0] _T_255; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [11:0] _T_256; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [11:0] _T_257; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [11:0] _T_258; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [11:0] _T_259; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [11:0] _T_260; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [11:0] _T_261; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [11:0] _T_262; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_263; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_264; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [51:0] _T_265; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [51:0] _T_266; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [51:0] _T_268; // @[Bitwise.scala 71:12]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [12:0] _T_269; // @[Cat.scala 29:58]
  wire [1:0] _T_271; // @[Cat.scala 29:58]
  wire [2:0] _T_273; // @[Cat.scala 29:58]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[55]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign _T_5 = ~io_in_sExp[11]; // @[primitives.scala 57:25]
  assign _T_7 = ~io_in_sExp[10]; // @[primitives.scala 57:25]
  assign _T_9 = ~io_in_sExp[9]; // @[primitives.scala 57:25]
  assign _T_11 = ~io_in_sExp[8]; // @[primitives.scala 57:25]
  assign _T_13 = ~io_in_sExp[7]; // @[primitives.scala 57:25]
  assign _T_15 = ~io_in_sExp[6]; // @[primitives.scala 57:25]
  assign _T_16 = ~io_in_sExp[5:0]; // @[primitives.scala 58:26]
  assign _T_17 = -65'sh10000000000000000 >>> _T_16; // @[primitives.scala 77:58]
  assign _T_23 = {{16'd0}, _T_17[44:29]}; // @[Bitwise.scala 102:31]
  assign _T_25 = {_T_17[28:13], 16'h0}; // @[Bitwise.scala 102:65]
  assign _T_27 = _T_25 & 32'hffff0000; // @[Bitwise.scala 102:75]
  assign _T_28 = _T_23 | _T_27; // @[Bitwise.scala 102:39]
  assign _GEN_0 = {{8'd0}, _T_28[31:8]}; // @[Bitwise.scala 102:31]
  assign _T_33 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 102:31]
  assign _T_35 = {_T_28[23:0], 8'h0}; // @[Bitwise.scala 102:65]
  assign _T_37 = _T_35 & 32'hff00ff00; // @[Bitwise.scala 102:75]
  assign _T_38 = _T_33 | _T_37; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{4'd0}, _T_38[31:4]}; // @[Bitwise.scala 102:31]
  assign _T_43 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 102:31]
  assign _T_45 = {_T_38[27:0], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_47 = _T_45 & 32'hf0f0f0f0; // @[Bitwise.scala 102:75]
  assign _T_48 = _T_43 | _T_47; // @[Bitwise.scala 102:39]
  assign _GEN_2 = {{2'd0}, _T_48[31:2]}; // @[Bitwise.scala 102:31]
  assign _T_53 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 102:31]
  assign _T_55 = {_T_48[29:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_57 = _T_55 & 32'hcccccccc; // @[Bitwise.scala 102:75]
  assign _T_58 = _T_53 | _T_57; // @[Bitwise.scala 102:39]
  assign _GEN_3 = {{1'd0}, _T_58[31:1]}; // @[Bitwise.scala 102:31]
  assign _T_63 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 102:31]
  assign _T_65 = {_T_58[30:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_67 = _T_65 & 32'haaaaaaaa; // @[Bitwise.scala 102:75]
  assign _T_68 = _T_63 | _T_67; // @[Bitwise.scala 102:39]
  assign _T_74 = {{8'd0}, _T_17[60:53]}; // @[Bitwise.scala 102:31]
  assign _T_76 = {_T_17[52:45], 8'h0}; // @[Bitwise.scala 102:65]
  assign _T_78 = _T_76 & 16'hff00; // @[Bitwise.scala 102:75]
  assign _T_79 = _T_74 | _T_78; // @[Bitwise.scala 102:39]
  assign _GEN_4 = {{4'd0}, _T_79[15:4]}; // @[Bitwise.scala 102:31]
  assign _T_84 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 102:31]
  assign _T_86 = {_T_79[11:0], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_88 = _T_86 & 16'hf0f0; // @[Bitwise.scala 102:75]
  assign _T_89 = _T_84 | _T_88; // @[Bitwise.scala 102:39]
  assign _GEN_5 = {{2'd0}, _T_89[15:2]}; // @[Bitwise.scala 102:31]
  assign _T_94 = _GEN_5 & 16'h3333; // @[Bitwise.scala 102:31]
  assign _T_96 = {_T_89[13:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_98 = _T_96 & 16'hcccc; // @[Bitwise.scala 102:75]
  assign _T_99 = _T_94 | _T_98; // @[Bitwise.scala 102:39]
  assign _GEN_6 = {{1'd0}, _T_99[15:1]}; // @[Bitwise.scala 102:31]
  assign _T_104 = _GEN_6 & 16'h5555; // @[Bitwise.scala 102:31]
  assign _T_106 = {_T_99[14:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_108 = _T_106 & 16'haaaa; // @[Bitwise.scala 102:75]
  assign _T_109 = _T_104 | _T_108; // @[Bitwise.scala 102:39]
  assign _T_118 = {_T_68,_T_109,_T_17[61],_T_17[62],_T_17[63]}; // @[Cat.scala 29:58]
  assign _T_120 = _T_15 ? 51'h0 : ~_T_118; // @[primitives.scala 74:21]
  assign _T_123 = _T_13 ? 51'h0 : _T_120[50:0]; // @[primitives.scala 74:21]
  assign _T_126 = _T_11 ? 51'h0 : _T_123[50:0]; // @[primitives.scala 74:21]
  assign _T_129 = _T_9 ? 51'h0 : _T_126[50:0]; // @[primitives.scala 74:21]
  assign _T_131 = {~_T_129,3'h7}; // @[Cat.scala 29:58]
  assign _T_147 = {_T_17[0],_T_17[1],_T_17[2]}; // @[Cat.scala 29:58]
  assign _T_148 = _T_15 ? _T_147 : 3'h0; // @[primitives.scala 61:24]
  assign _T_149 = _T_13 ? _T_148 : 3'h0; // @[primitives.scala 61:24]
  assign _T_150 = _T_11 ? _T_149 : 3'h0; // @[primitives.scala 61:24]
  assign _T_151 = _T_9 ? _T_150 : 3'h0; // @[primitives.scala 61:24]
  assign _T_152 = _T_7 ? _T_131 : {{51'd0}, _T_151}; // @[primitives.scala 66:24]
  assign _T_153 = _T_5 ? _T_152 : 54'h0; // @[primitives.scala 61:24]
  assign _GEN_7 = {{53'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_154 = _T_153 | _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_155 = {_T_154,2'h3}; // @[Cat.scala 29:58]
  assign _T_157 = {1'h0,_T_155[55:1]}; // @[Cat.scala 29:58]
  assign _T_159 = ~_T_157 & _T_155; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_160 = io_in_sig & _T_159; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_161 = _T_160 != 56'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_162 = io_in_sig & _T_157; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_163 = _T_162 != 56'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_164 = _T_161 | _T_163; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_165 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_166 = _T_165 & _T_161; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_167 = roundMagUp & _T_164; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_168 = _T_166 | _T_167; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_169 = io_in_sig | _T_155; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_171 = _T_169[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_172 = roundingMode_near_even & _T_161; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_174 = _T_172 & ~_T_163; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_176 = _T_174 ? _T_155[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_178 = _T_171 & ~_T_176; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_180 = io_in_sig & ~_T_155; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_182 = roundingMode_odd & _T_164; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_184 = _T_182 ? _T_159[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_8 = {{1'd0}, _T_180[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_185 = _GEN_8 | _T_184; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_186 = _T_168 ? _T_178 : _T_185; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_188 = {1'b0,$signed(_T_186[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_9 = {{10{_T_188[2]}},_T_188}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_189 = $signed(io_in_sExp) + $signed(_GEN_9); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_189[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? _T_186[52:1] : _T_186[51:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _T_194 = _T_189[13:10]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_194) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_189) < 14'sh3ce; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_199 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _T_201 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _T_203 = io_in_sig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_204 = _T_201 | _T_203; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _T_206 = _T_165 & _T_199; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_207 = roundMagUp & _T_204; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_208 = _T_206 | _T_207; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_211 = doShiftSigDown1 ? _T_186[54] : _T_186[53]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _T_212 = io_in_sExp[12:11]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_213 = $signed(_T_212) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_214 = _T_164 & _T_213; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_217 = doShiftSigDown1 ? _T_155[3] : _T_155[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _T_218 = _T_214 & _T_217; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_222 = doShiftSigDown1 ? _T_155[4] : _T_155[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _T_224 = io_detectTininess & ~_T_222; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_225 = _T_224 & _T_211; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_226 = _T_225 & _T_161; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_227 = _T_226 & _T_208; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_229 = _T_218 & ~_T_227; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_229; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_164; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign _T_234 = ~isNaNOut & ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_234 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_236 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_236; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_165 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_238 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_239 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_238 & _T_239; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_241 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = io_in_isInf | _T_241; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_242 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_243 = _T_242 ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_245 = common_expOut & ~_T_243; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_247 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_249 = _T_245 & ~_T_247; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_250 = pegMaxFiniteMagOut ? 12'h400 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_252 = _T_249 & ~_T_250; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_253 = notNaN_isInfOut ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_255 = _T_252 & ~_T_253; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_256 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_257 = _T_255 | _T_256; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_258 = pegMaxFiniteMagOut ? 12'hbff : 12'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_259 = _T_257 | _T_258; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_260 = notNaN_isInfOut ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_261 = _T_259 | _T_260; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_262 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_261 | _T_262; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_263 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_264 = _T_263 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_265 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_266 = _T_264 ? _T_265 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_268 = pegMaxFiniteMagOut ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 71:12]
  assign fractOut = _T_266 | _T_268; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_269 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_271 = {underflow,inexact}; // @[Cat.scala 29:58]
  assign _T_273 = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_269,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_273,_T_271}; // @[RoundAnyRawFNToRecFN.scala 285:23]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [12:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [55:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
endmodule
module MulAddRecFN(
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire [64:0] mulAddRecFNToRaw_preMul_io_a; // @[MulAddRecFN.scala 318:15]
  wire [64:0] mulAddRecFNToRaw_preMul_io_b; // @[MulAddRecFN.scala 318:15]
  wire [64:0] mulAddRecFNToRaw_preMul_io_c; // @[MulAddRecFN.scala 318:15]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[MulAddRecFN.scala 318:15]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 318:15]
  wire [105:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 318:15]
  wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 318:15]
  wire [5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 318:15]
  wire [54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 320:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 320:15]
  wire [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 320:15]
  wire [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[MulAddRecFN.scala 320:15]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 320:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 320:15]
  wire [55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 320:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulAddRecFN.scala 340:15]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[MulAddRecFN.scala 340:15]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[MulAddRecFN.scala 340:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[MulAddRecFN.scala 340:15]
  wire [64:0] roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 340:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[MulAddRecFN.scala 340:15]
  wire [105:0] _T; // @[MulAddRecFN.scala 328:45]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[MulAddRecFN.scala 318:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[MulAddRecFN.scala 320:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[MulAddRecFN.scala 340:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags)
  );
  assign _T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 328:45]
  assign io_out = roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 346:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[MulAddRecFN.scala 347:23]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[MulAddRecFN.scala 323:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[MulAddRecFN.scala 324:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[MulAddRecFN.scala 325:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 334:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = io_roundingMode; // @[MulAddRecFN.scala 335:46]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 341:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_roundingMode = io_roundingMode; // @[MulAddRecFN.scala 344:39]
  assign roundRawFNToRecFN_io_detectTininess = io_detectTininess; // @[MulAddRecFN.scala 345:41]
endmodule
module ValExec_MulAddRecF64_mul(
  input         clock,
  input         reset,
  input  [63:0] io_a,
  input  [63:0] io_b,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [63:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [64:0] io_expected_recOut,
  output [64:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [64:0] mulAddRecFN_io_a; // @[ValExec_MulAddRecFN.scala 158:29]
  wire [64:0] mulAddRecFN_io_b; // @[ValExec_MulAddRecFN.scala 158:29]
  wire [64:0] mulAddRecFN_io_c; // @[ValExec_MulAddRecFN.scala 158:29]
  wire [2:0] mulAddRecFN_io_roundingMode; // @[ValExec_MulAddRecFN.scala 158:29]
  wire  mulAddRecFN_io_detectTininess; // @[ValExec_MulAddRecFN.scala 158:29]
  wire [64:0] mulAddRecFN_io_out; // @[ValExec_MulAddRecFN.scala 158:29]
  wire [4:0] mulAddRecFN_io_exceptionFlags; // @[ValExec_MulAddRecFN.scala 158:29]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_57; // @[Mux.scala 47:69]
  wire [5:0] _T_58; // @[Mux.scala 47:69]
  wire [5:0] _T_59; // @[Mux.scala 47:69]
  wire [5:0] _T_60; // @[Mux.scala 47:69]
  wire [5:0] _T_61; // @[Mux.scala 47:69]
  wire [5:0] _T_62; // @[Mux.scala 47:69]
  wire [5:0] _T_63; // @[Mux.scala 47:69]
  wire [5:0] _T_64; // @[Mux.scala 47:69]
  wire [5:0] _T_65; // @[Mux.scala 47:69]
  wire [5:0] _T_66; // @[Mux.scala 47:69]
  wire [5:0] _T_67; // @[Mux.scala 47:69]
  wire [5:0] _T_68; // @[Mux.scala 47:69]
  wire [5:0] _T_69; // @[Mux.scala 47:69]
  wire [5:0] _T_70; // @[Mux.scala 47:69]
  wire [5:0] _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [114:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_108; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_110; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_111; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_112; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_113; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_114; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_116; // @[rawFloatFromFN.scala 59:15]
  wire  _T_117; // @[rawFloatFromFN.scala 62:34]
  wire  _T_119; // @[rawFloatFromFN.scala 63:62]
  wire  _T_122; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_125; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_127; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_129; // @[Cat.scala 29:58]
  wire [2:0] _T_131; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_133; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_136; // @[Cat.scala 29:58]
  wire [3:0] _T_137; // @[Cat.scala 29:58]
  wire  _T_142; // @[rawFloatFromFN.scala 50:34]
  wire  _T_143; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_196; // @[Mux.scala 47:69]
  wire [5:0] _T_197; // @[Mux.scala 47:69]
  wire [5:0] _T_198; // @[Mux.scala 47:69]
  wire [5:0] _T_199; // @[Mux.scala 47:69]
  wire [5:0] _T_200; // @[Mux.scala 47:69]
  wire [5:0] _T_201; // @[Mux.scala 47:69]
  wire [5:0] _T_202; // @[Mux.scala 47:69]
  wire [5:0] _T_203; // @[Mux.scala 47:69]
  wire [5:0] _T_204; // @[Mux.scala 47:69]
  wire [5:0] _T_205; // @[Mux.scala 47:69]
  wire [5:0] _T_206; // @[Mux.scala 47:69]
  wire [5:0] _T_207; // @[Mux.scala 47:69]
  wire [5:0] _T_208; // @[Mux.scala 47:69]
  wire [5:0] _T_209; // @[Mux.scala 47:69]
  wire [5:0] _T_210; // @[Mux.scala 47:69]
  wire [5:0] _T_211; // @[Mux.scala 47:69]
  wire [5:0] _T_212; // @[Mux.scala 47:69]
  wire [5:0] _T_213; // @[Mux.scala 47:69]
  wire [5:0] _T_214; // @[Mux.scala 47:69]
  wire [5:0] _T_215; // @[Mux.scala 47:69]
  wire [5:0] _T_216; // @[Mux.scala 47:69]
  wire [5:0] _T_217; // @[Mux.scala 47:69]
  wire [5:0] _T_218; // @[Mux.scala 47:69]
  wire [5:0] _T_219; // @[Mux.scala 47:69]
  wire [5:0] _T_220; // @[Mux.scala 47:69]
  wire [5:0] _T_221; // @[Mux.scala 47:69]
  wire [5:0] _T_222; // @[Mux.scala 47:69]
  wire [5:0] _T_223; // @[Mux.scala 47:69]
  wire [5:0] _T_224; // @[Mux.scala 47:69]
  wire [5:0] _T_225; // @[Mux.scala 47:69]
  wire [5:0] _T_226; // @[Mux.scala 47:69]
  wire [5:0] _T_227; // @[Mux.scala 47:69]
  wire [5:0] _T_228; // @[Mux.scala 47:69]
  wire [5:0] _T_229; // @[Mux.scala 47:69]
  wire [5:0] _T_230; // @[Mux.scala 47:69]
  wire [5:0] _T_231; // @[Mux.scala 47:69]
  wire [5:0] _T_232; // @[Mux.scala 47:69]
  wire [5:0] _T_233; // @[Mux.scala 47:69]
  wire [5:0] _T_234; // @[Mux.scala 47:69]
  wire [5:0] _T_235; // @[Mux.scala 47:69]
  wire [5:0] _T_236; // @[Mux.scala 47:69]
  wire [5:0] _T_237; // @[Mux.scala 47:69]
  wire [5:0] _T_238; // @[Mux.scala 47:69]
  wire [5:0] _T_239; // @[Mux.scala 47:69]
  wire [5:0] _T_240; // @[Mux.scala 47:69]
  wire [5:0] _T_241; // @[Mux.scala 47:69]
  wire [5:0] _T_242; // @[Mux.scala 47:69]
  wire [5:0] _T_243; // @[Mux.scala 47:69]
  wire [5:0] _T_244; // @[Mux.scala 47:69]
  wire [5:0] _T_245; // @[Mux.scala 47:69]
  wire [5:0] _T_246; // @[Mux.scala 47:69]
  wire [114:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_247; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_249; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_250; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_251; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_252; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_253; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_255; // @[rawFloatFromFN.scala 59:15]
  wire  _T_256; // @[rawFloatFromFN.scala 62:34]
  wire  _T_258; // @[rawFloatFromFN.scala 63:62]
  wire  _T_261; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_264; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_266; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_268; // @[Cat.scala 29:58]
  wire [2:0] _T_270; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_272; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_275; // @[Cat.scala 29:58]
  wire [3:0] _T_276; // @[Cat.scala 29:58]
  wire [63:0] _T_278; // @[ValExec_MulAddRecFN.scala 163:16]
  wire [63:0] _T_279; // @[ValExec_MulAddRecFN.scala 163:24]
  wire  _T_284; // @[rawFloatFromFN.scala 50:34]
  wire  _T_285; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_338; // @[Mux.scala 47:69]
  wire [5:0] _T_339; // @[Mux.scala 47:69]
  wire [5:0] _T_340; // @[Mux.scala 47:69]
  wire [5:0] _T_341; // @[Mux.scala 47:69]
  wire [5:0] _T_342; // @[Mux.scala 47:69]
  wire [5:0] _T_343; // @[Mux.scala 47:69]
  wire [5:0] _T_344; // @[Mux.scala 47:69]
  wire [5:0] _T_345; // @[Mux.scala 47:69]
  wire [5:0] _T_346; // @[Mux.scala 47:69]
  wire [5:0] _T_347; // @[Mux.scala 47:69]
  wire [5:0] _T_348; // @[Mux.scala 47:69]
  wire [5:0] _T_349; // @[Mux.scala 47:69]
  wire [5:0] _T_350; // @[Mux.scala 47:69]
  wire [5:0] _T_351; // @[Mux.scala 47:69]
  wire [5:0] _T_352; // @[Mux.scala 47:69]
  wire [5:0] _T_353; // @[Mux.scala 47:69]
  wire [5:0] _T_354; // @[Mux.scala 47:69]
  wire [5:0] _T_355; // @[Mux.scala 47:69]
  wire [5:0] _T_356; // @[Mux.scala 47:69]
  wire [5:0] _T_357; // @[Mux.scala 47:69]
  wire [5:0] _T_358; // @[Mux.scala 47:69]
  wire [5:0] _T_359; // @[Mux.scala 47:69]
  wire [5:0] _T_360; // @[Mux.scala 47:69]
  wire [5:0] _T_361; // @[Mux.scala 47:69]
  wire [5:0] _T_362; // @[Mux.scala 47:69]
  wire [5:0] _T_363; // @[Mux.scala 47:69]
  wire [5:0] _T_364; // @[Mux.scala 47:69]
  wire [5:0] _T_365; // @[Mux.scala 47:69]
  wire [5:0] _T_366; // @[Mux.scala 47:69]
  wire [5:0] _T_367; // @[Mux.scala 47:69]
  wire [5:0] _T_368; // @[Mux.scala 47:69]
  wire [5:0] _T_369; // @[Mux.scala 47:69]
  wire [5:0] _T_370; // @[Mux.scala 47:69]
  wire [5:0] _T_371; // @[Mux.scala 47:69]
  wire [5:0] _T_372; // @[Mux.scala 47:69]
  wire [5:0] _T_373; // @[Mux.scala 47:69]
  wire [5:0] _T_374; // @[Mux.scala 47:69]
  wire [5:0] _T_375; // @[Mux.scala 47:69]
  wire [5:0] _T_376; // @[Mux.scala 47:69]
  wire [5:0] _T_377; // @[Mux.scala 47:69]
  wire [5:0] _T_378; // @[Mux.scala 47:69]
  wire [5:0] _T_379; // @[Mux.scala 47:69]
  wire [5:0] _T_380; // @[Mux.scala 47:69]
  wire [5:0] _T_381; // @[Mux.scala 47:69]
  wire [5:0] _T_382; // @[Mux.scala 47:69]
  wire [5:0] _T_383; // @[Mux.scala 47:69]
  wire [5:0] _T_384; // @[Mux.scala 47:69]
  wire [5:0] _T_385; // @[Mux.scala 47:69]
  wire [5:0] _T_386; // @[Mux.scala 47:69]
  wire [5:0] _T_387; // @[Mux.scala 47:69]
  wire [5:0] _T_388; // @[Mux.scala 47:69]
  wire [114:0] _GEN_10; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_389; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_391; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_11; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_392; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_393; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_394; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_12; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_395; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_13; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_397; // @[rawFloatFromFN.scala 59:15]
  wire  _T_398; // @[rawFloatFromFN.scala 62:34]
  wire  _T_400; // @[rawFloatFromFN.scala 63:62]
  wire  _T_403; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_406; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_408; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_410; // @[Cat.scala 29:58]
  wire [2:0] _T_412; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_14; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_414; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_417; // @[Cat.scala 29:58]
  wire [3:0] _T_418; // @[Cat.scala 29:58]
  wire  _T_423; // @[tests.scala 48:26]
  wire  _T_425; // @[tests.scala 48:55]
  wire  _T_426; // @[tests.scala 48:39]
  wire  _T_427; // @[tests.scala 49:20]
  wire  _T_430; // @[tests.scala 49:54]
  wire  _T_431; // @[tests.scala 49:31]
  wire  _T_433; // @[tests.scala 50:30]
  wire  _T_435; // @[tests.scala 50:66]
  wire  _T_436; // @[tests.scala 50:16]
  wire  _T_437; // @[tests.scala 48:12]
  wire  _T_438; // @[ValExec_MulAddRecFN.scala 175:35]
  MulAddRecFN mulAddRecFN ( // @[ValExec_MulAddRecFN.scala 158:29]
    .io_a(mulAddRecFN_io_a),
    .io_b(mulAddRecFN_io_b),
    .io_c(mulAddRecFN_io_c),
    .io_roundingMode(mulAddRecFN_io_roundingMode),
    .io_detectTininess(mulAddRecFN_io_detectTininess),
    .io_out(mulAddRecFN_io_out),
    .io_exceptionFlags(mulAddRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_a[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_a[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_57 = io_a[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_58 = io_a[2] ? 6'h31 : _T_57; // @[Mux.scala 47:69]
  assign _T_59 = io_a[3] ? 6'h30 : _T_58; // @[Mux.scala 47:69]
  assign _T_60 = io_a[4] ? 6'h2f : _T_59; // @[Mux.scala 47:69]
  assign _T_61 = io_a[5] ? 6'h2e : _T_60; // @[Mux.scala 47:69]
  assign _T_62 = io_a[6] ? 6'h2d : _T_61; // @[Mux.scala 47:69]
  assign _T_63 = io_a[7] ? 6'h2c : _T_62; // @[Mux.scala 47:69]
  assign _T_64 = io_a[8] ? 6'h2b : _T_63; // @[Mux.scala 47:69]
  assign _T_65 = io_a[9] ? 6'h2a : _T_64; // @[Mux.scala 47:69]
  assign _T_66 = io_a[10] ? 6'h29 : _T_65; // @[Mux.scala 47:69]
  assign _T_67 = io_a[11] ? 6'h28 : _T_66; // @[Mux.scala 47:69]
  assign _T_68 = io_a[12] ? 6'h27 : _T_67; // @[Mux.scala 47:69]
  assign _T_69 = io_a[13] ? 6'h26 : _T_68; // @[Mux.scala 47:69]
  assign _T_70 = io_a[14] ? 6'h25 : _T_69; // @[Mux.scala 47:69]
  assign _T_71 = io_a[15] ? 6'h24 : _T_70; // @[Mux.scala 47:69]
  assign _T_72 = io_a[16] ? 6'h23 : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = io_a[17] ? 6'h22 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = io_a[18] ? 6'h21 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = io_a[19] ? 6'h20 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = io_a[20] ? 6'h1f : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = io_a[21] ? 6'h1e : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = io_a[22] ? 6'h1d : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = io_a[23] ? 6'h1c : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = io_a[24] ? 6'h1b : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = io_a[25] ? 6'h1a : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = io_a[26] ? 6'h19 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = io_a[27] ? 6'h18 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = io_a[28] ? 6'h17 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = io_a[29] ? 6'h16 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = io_a[30] ? 6'h15 : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = io_a[31] ? 6'h14 : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = io_a[32] ? 6'h13 : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = io_a[33] ? 6'h12 : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = io_a[34] ? 6'h11 : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = io_a[35] ? 6'h10 : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = io_a[36] ? 6'hf : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = io_a[37] ? 6'he : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = io_a[38] ? 6'hd : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = io_a[39] ? 6'hc : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = io_a[40] ? 6'hb : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = io_a[41] ? 6'ha : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = io_a[42] ? 6'h9 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = io_a[43] ? 6'h8 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = io_a[44] ? 6'h7 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = io_a[45] ? 6'h6 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = io_a[46] ? 6'h5 : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = io_a[47] ? 6'h4 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = io_a[48] ? 6'h3 : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = io_a[49] ? 6'h2 : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = io_a[50] ? 6'h1 : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = io_a[51] ? 6'h0 : _T_106; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, io_a[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_108 = _GEN_0 << _T_107; // @[rawFloatFromFN.scala 54:36]
  assign _T_110 = {_T_108[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{6'd0}, _T_107}; // @[rawFloatFromFN.scala 57:26]
  assign _T_111 = _GEN_1 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_112 = _T_3 ? _T_111 : {{1'd0}, io_a[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_113 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{9'd0}, _T_113}; // @[rawFloatFromFN.scala 60:22]
  assign _T_114 = 11'h400 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_114}; // @[rawFloatFromFN.scala 59:15]
  assign _T_116 = _T_112 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_117 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_119 = _T_116[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_122 = _T_119 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_125 = {1'b0,$signed(_T_116)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_127 = _T_3 ? _T_110 : io_a[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_129 = {1'h0,~_T_117,_T_127}; // @[Cat.scala 29:58]
  assign _T_131 = _T_117 ? 3'h0 : _T_125[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_122}; // @[recFNFromFN.scala 48:79]
  assign _T_133 = _T_131 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_136 = {_T_125[8:0],_T_129[51:0]}; // @[Cat.scala 29:58]
  assign _T_137 = {io_a[63],_T_133}; // @[Cat.scala 29:58]
  assign _T_142 = io_b[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_143 = io_b[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_196 = io_b[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_197 = io_b[2] ? 6'h31 : _T_196; // @[Mux.scala 47:69]
  assign _T_198 = io_b[3] ? 6'h30 : _T_197; // @[Mux.scala 47:69]
  assign _T_199 = io_b[4] ? 6'h2f : _T_198; // @[Mux.scala 47:69]
  assign _T_200 = io_b[5] ? 6'h2e : _T_199; // @[Mux.scala 47:69]
  assign _T_201 = io_b[6] ? 6'h2d : _T_200; // @[Mux.scala 47:69]
  assign _T_202 = io_b[7] ? 6'h2c : _T_201; // @[Mux.scala 47:69]
  assign _T_203 = io_b[8] ? 6'h2b : _T_202; // @[Mux.scala 47:69]
  assign _T_204 = io_b[9] ? 6'h2a : _T_203; // @[Mux.scala 47:69]
  assign _T_205 = io_b[10] ? 6'h29 : _T_204; // @[Mux.scala 47:69]
  assign _T_206 = io_b[11] ? 6'h28 : _T_205; // @[Mux.scala 47:69]
  assign _T_207 = io_b[12] ? 6'h27 : _T_206; // @[Mux.scala 47:69]
  assign _T_208 = io_b[13] ? 6'h26 : _T_207; // @[Mux.scala 47:69]
  assign _T_209 = io_b[14] ? 6'h25 : _T_208; // @[Mux.scala 47:69]
  assign _T_210 = io_b[15] ? 6'h24 : _T_209; // @[Mux.scala 47:69]
  assign _T_211 = io_b[16] ? 6'h23 : _T_210; // @[Mux.scala 47:69]
  assign _T_212 = io_b[17] ? 6'h22 : _T_211; // @[Mux.scala 47:69]
  assign _T_213 = io_b[18] ? 6'h21 : _T_212; // @[Mux.scala 47:69]
  assign _T_214 = io_b[19] ? 6'h20 : _T_213; // @[Mux.scala 47:69]
  assign _T_215 = io_b[20] ? 6'h1f : _T_214; // @[Mux.scala 47:69]
  assign _T_216 = io_b[21] ? 6'h1e : _T_215; // @[Mux.scala 47:69]
  assign _T_217 = io_b[22] ? 6'h1d : _T_216; // @[Mux.scala 47:69]
  assign _T_218 = io_b[23] ? 6'h1c : _T_217; // @[Mux.scala 47:69]
  assign _T_219 = io_b[24] ? 6'h1b : _T_218; // @[Mux.scala 47:69]
  assign _T_220 = io_b[25] ? 6'h1a : _T_219; // @[Mux.scala 47:69]
  assign _T_221 = io_b[26] ? 6'h19 : _T_220; // @[Mux.scala 47:69]
  assign _T_222 = io_b[27] ? 6'h18 : _T_221; // @[Mux.scala 47:69]
  assign _T_223 = io_b[28] ? 6'h17 : _T_222; // @[Mux.scala 47:69]
  assign _T_224 = io_b[29] ? 6'h16 : _T_223; // @[Mux.scala 47:69]
  assign _T_225 = io_b[30] ? 6'h15 : _T_224; // @[Mux.scala 47:69]
  assign _T_226 = io_b[31] ? 6'h14 : _T_225; // @[Mux.scala 47:69]
  assign _T_227 = io_b[32] ? 6'h13 : _T_226; // @[Mux.scala 47:69]
  assign _T_228 = io_b[33] ? 6'h12 : _T_227; // @[Mux.scala 47:69]
  assign _T_229 = io_b[34] ? 6'h11 : _T_228; // @[Mux.scala 47:69]
  assign _T_230 = io_b[35] ? 6'h10 : _T_229; // @[Mux.scala 47:69]
  assign _T_231 = io_b[36] ? 6'hf : _T_230; // @[Mux.scala 47:69]
  assign _T_232 = io_b[37] ? 6'he : _T_231; // @[Mux.scala 47:69]
  assign _T_233 = io_b[38] ? 6'hd : _T_232; // @[Mux.scala 47:69]
  assign _T_234 = io_b[39] ? 6'hc : _T_233; // @[Mux.scala 47:69]
  assign _T_235 = io_b[40] ? 6'hb : _T_234; // @[Mux.scala 47:69]
  assign _T_236 = io_b[41] ? 6'ha : _T_235; // @[Mux.scala 47:69]
  assign _T_237 = io_b[42] ? 6'h9 : _T_236; // @[Mux.scala 47:69]
  assign _T_238 = io_b[43] ? 6'h8 : _T_237; // @[Mux.scala 47:69]
  assign _T_239 = io_b[44] ? 6'h7 : _T_238; // @[Mux.scala 47:69]
  assign _T_240 = io_b[45] ? 6'h6 : _T_239; // @[Mux.scala 47:69]
  assign _T_241 = io_b[46] ? 6'h5 : _T_240; // @[Mux.scala 47:69]
  assign _T_242 = io_b[47] ? 6'h4 : _T_241; // @[Mux.scala 47:69]
  assign _T_243 = io_b[48] ? 6'h3 : _T_242; // @[Mux.scala 47:69]
  assign _T_244 = io_b[49] ? 6'h2 : _T_243; // @[Mux.scala 47:69]
  assign _T_245 = io_b[50] ? 6'h1 : _T_244; // @[Mux.scala 47:69]
  assign _T_246 = io_b[51] ? 6'h0 : _T_245; // @[Mux.scala 47:69]
  assign _GEN_5 = {{63'd0}, io_b[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_247 = _GEN_5 << _T_246; // @[rawFloatFromFN.scala 54:36]
  assign _T_249 = {_T_247[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{6'd0}, _T_246}; // @[rawFloatFromFN.scala 57:26]
  assign _T_250 = _GEN_6 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_251 = _T_142 ? _T_250 : {{1'd0}, io_b[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_252 = _T_142 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{9'd0}, _T_252}; // @[rawFloatFromFN.scala 60:22]
  assign _T_253 = 11'h400 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_253}; // @[rawFloatFromFN.scala 59:15]
  assign _T_255 = _T_251 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_256 = _T_142 & _T_143; // @[rawFloatFromFN.scala 62:34]
  assign _T_258 = _T_255[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_261 = _T_258 & ~_T_143; // @[rawFloatFromFN.scala 66:33]
  assign _T_264 = {1'b0,$signed(_T_255)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_266 = _T_142 ? _T_249 : io_b[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_268 = {1'h0,~_T_256,_T_266}; // @[Cat.scala 29:58]
  assign _T_270 = _T_256 ? 3'h0 : _T_264[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_261}; // @[recFNFromFN.scala 48:79]
  assign _T_272 = _T_270 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_275 = {_T_264[8:0],_T_268[51:0]}; // @[Cat.scala 29:58]
  assign _T_276 = {io_b[63],_T_272}; // @[Cat.scala 29:58]
  assign _T_278 = io_a ^ io_b; // @[ValExec_MulAddRecFN.scala 163:16]
  assign _T_279 = _T_278 & 64'h8000000000000000; // @[ValExec_MulAddRecFN.scala 163:24]
  assign _T_284 = io_expected_out[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_285 = io_expected_out[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_338 = io_expected_out[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_339 = io_expected_out[2] ? 6'h31 : _T_338; // @[Mux.scala 47:69]
  assign _T_340 = io_expected_out[3] ? 6'h30 : _T_339; // @[Mux.scala 47:69]
  assign _T_341 = io_expected_out[4] ? 6'h2f : _T_340; // @[Mux.scala 47:69]
  assign _T_342 = io_expected_out[5] ? 6'h2e : _T_341; // @[Mux.scala 47:69]
  assign _T_343 = io_expected_out[6] ? 6'h2d : _T_342; // @[Mux.scala 47:69]
  assign _T_344 = io_expected_out[7] ? 6'h2c : _T_343; // @[Mux.scala 47:69]
  assign _T_345 = io_expected_out[8] ? 6'h2b : _T_344; // @[Mux.scala 47:69]
  assign _T_346 = io_expected_out[9] ? 6'h2a : _T_345; // @[Mux.scala 47:69]
  assign _T_347 = io_expected_out[10] ? 6'h29 : _T_346; // @[Mux.scala 47:69]
  assign _T_348 = io_expected_out[11] ? 6'h28 : _T_347; // @[Mux.scala 47:69]
  assign _T_349 = io_expected_out[12] ? 6'h27 : _T_348; // @[Mux.scala 47:69]
  assign _T_350 = io_expected_out[13] ? 6'h26 : _T_349; // @[Mux.scala 47:69]
  assign _T_351 = io_expected_out[14] ? 6'h25 : _T_350; // @[Mux.scala 47:69]
  assign _T_352 = io_expected_out[15] ? 6'h24 : _T_351; // @[Mux.scala 47:69]
  assign _T_353 = io_expected_out[16] ? 6'h23 : _T_352; // @[Mux.scala 47:69]
  assign _T_354 = io_expected_out[17] ? 6'h22 : _T_353; // @[Mux.scala 47:69]
  assign _T_355 = io_expected_out[18] ? 6'h21 : _T_354; // @[Mux.scala 47:69]
  assign _T_356 = io_expected_out[19] ? 6'h20 : _T_355; // @[Mux.scala 47:69]
  assign _T_357 = io_expected_out[20] ? 6'h1f : _T_356; // @[Mux.scala 47:69]
  assign _T_358 = io_expected_out[21] ? 6'h1e : _T_357; // @[Mux.scala 47:69]
  assign _T_359 = io_expected_out[22] ? 6'h1d : _T_358; // @[Mux.scala 47:69]
  assign _T_360 = io_expected_out[23] ? 6'h1c : _T_359; // @[Mux.scala 47:69]
  assign _T_361 = io_expected_out[24] ? 6'h1b : _T_360; // @[Mux.scala 47:69]
  assign _T_362 = io_expected_out[25] ? 6'h1a : _T_361; // @[Mux.scala 47:69]
  assign _T_363 = io_expected_out[26] ? 6'h19 : _T_362; // @[Mux.scala 47:69]
  assign _T_364 = io_expected_out[27] ? 6'h18 : _T_363; // @[Mux.scala 47:69]
  assign _T_365 = io_expected_out[28] ? 6'h17 : _T_364; // @[Mux.scala 47:69]
  assign _T_366 = io_expected_out[29] ? 6'h16 : _T_365; // @[Mux.scala 47:69]
  assign _T_367 = io_expected_out[30] ? 6'h15 : _T_366; // @[Mux.scala 47:69]
  assign _T_368 = io_expected_out[31] ? 6'h14 : _T_367; // @[Mux.scala 47:69]
  assign _T_369 = io_expected_out[32] ? 6'h13 : _T_368; // @[Mux.scala 47:69]
  assign _T_370 = io_expected_out[33] ? 6'h12 : _T_369; // @[Mux.scala 47:69]
  assign _T_371 = io_expected_out[34] ? 6'h11 : _T_370; // @[Mux.scala 47:69]
  assign _T_372 = io_expected_out[35] ? 6'h10 : _T_371; // @[Mux.scala 47:69]
  assign _T_373 = io_expected_out[36] ? 6'hf : _T_372; // @[Mux.scala 47:69]
  assign _T_374 = io_expected_out[37] ? 6'he : _T_373; // @[Mux.scala 47:69]
  assign _T_375 = io_expected_out[38] ? 6'hd : _T_374; // @[Mux.scala 47:69]
  assign _T_376 = io_expected_out[39] ? 6'hc : _T_375; // @[Mux.scala 47:69]
  assign _T_377 = io_expected_out[40] ? 6'hb : _T_376; // @[Mux.scala 47:69]
  assign _T_378 = io_expected_out[41] ? 6'ha : _T_377; // @[Mux.scala 47:69]
  assign _T_379 = io_expected_out[42] ? 6'h9 : _T_378; // @[Mux.scala 47:69]
  assign _T_380 = io_expected_out[43] ? 6'h8 : _T_379; // @[Mux.scala 47:69]
  assign _T_381 = io_expected_out[44] ? 6'h7 : _T_380; // @[Mux.scala 47:69]
  assign _T_382 = io_expected_out[45] ? 6'h6 : _T_381; // @[Mux.scala 47:69]
  assign _T_383 = io_expected_out[46] ? 6'h5 : _T_382; // @[Mux.scala 47:69]
  assign _T_384 = io_expected_out[47] ? 6'h4 : _T_383; // @[Mux.scala 47:69]
  assign _T_385 = io_expected_out[48] ? 6'h3 : _T_384; // @[Mux.scala 47:69]
  assign _T_386 = io_expected_out[49] ? 6'h2 : _T_385; // @[Mux.scala 47:69]
  assign _T_387 = io_expected_out[50] ? 6'h1 : _T_386; // @[Mux.scala 47:69]
  assign _T_388 = io_expected_out[51] ? 6'h0 : _T_387; // @[Mux.scala 47:69]
  assign _GEN_10 = {{63'd0}, io_expected_out[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_389 = _GEN_10 << _T_388; // @[rawFloatFromFN.scala 54:36]
  assign _T_391 = {_T_389[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_11 = {{6'd0}, _T_388}; // @[rawFloatFromFN.scala 57:26]
  assign _T_392 = _GEN_11 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_393 = _T_284 ? _T_392 : {{1'd0}, io_expected_out[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_394 = _T_284 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_12 = {{9'd0}, _T_394}; // @[rawFloatFromFN.scala 60:22]
  assign _T_395 = 11'h400 | _GEN_12; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_13 = {{1'd0}, _T_395}; // @[rawFloatFromFN.scala 59:15]
  assign _T_397 = _T_393 + _GEN_13; // @[rawFloatFromFN.scala 59:15]
  assign _T_398 = _T_284 & _T_285; // @[rawFloatFromFN.scala 62:34]
  assign _T_400 = _T_397[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_403 = _T_400 & ~_T_285; // @[rawFloatFromFN.scala 66:33]
  assign _T_406 = {1'b0,$signed(_T_397)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_408 = _T_284 ? _T_391 : io_expected_out[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_410 = {1'h0,~_T_398,_T_408}; // @[Cat.scala 29:58]
  assign _T_412 = _T_398 ? 3'h0 : _T_406[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_14 = {{2'd0}, _T_403}; // @[recFNFromFN.scala 48:79]
  assign _T_414 = _T_412 | _GEN_14; // @[recFNFromFN.scala 48:79]
  assign _T_417 = {_T_406[8:0],_T_410[51:0]}; // @[Cat.scala 29:58]
  assign _T_418 = {io_expected_out[63],_T_414}; // @[Cat.scala 29:58]
  assign _T_423 = io_actual_out[63:61] == 3'h0; // @[tests.scala 48:26]
  assign _T_425 = io_actual_out[63:61] == 3'h7; // @[tests.scala 48:55]
  assign _T_426 = _T_423 | _T_425; // @[tests.scala 48:39]
  assign _T_427 = io_actual_out[64:61] == io_expected_recOut[64:61]; // @[tests.scala 49:20]
  assign _T_430 = io_actual_out[51:0] == io_expected_recOut[51:0]; // @[tests.scala 49:54]
  assign _T_431 = _T_427 & _T_430; // @[tests.scala 49:31]
  assign _T_433 = io_actual_out[63:61] == 3'h6; // @[tests.scala 50:30]
  assign _T_435 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_436 = _T_433 ? _T_427 : _T_435; // @[tests.scala 50:16]
  assign _T_437 = _T_426 ? _T_431 : _T_436; // @[tests.scala 48:12]
  assign _T_438 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_MulAddRecFN.scala 175:35]
  assign io_expected_recOut = {_T_418,_T_417}; // @[ValExec_MulAddRecFN.scala 167:24]
  assign io_actual_out = mulAddRecFN_io_out; // @[ValExec_MulAddRecFN.scala 169:19]
  assign io_actual_exceptionFlags = mulAddRecFN_io_exceptionFlags; // @[ValExec_MulAddRecFN.scala 170:30]
  assign io_check = 1'h1; // @[ValExec_MulAddRecFN.scala 172:14]
  assign io_pass = _T_437 & _T_438; // @[ValExec_MulAddRecFN.scala 173:13]
  assign mulAddRecFN_io_a = {_T_137,_T_136}; // @[ValExec_MulAddRecFN.scala 160:22]
  assign mulAddRecFN_io_b = {_T_276,_T_275}; // @[ValExec_MulAddRecFN.scala 161:22]
  assign mulAddRecFN_io_c = {_T_279, 1'h0}; // @[ValExec_MulAddRecFN.scala 162:22]
  assign mulAddRecFN_io_roundingMode = io_roundingMode; // @[ValExec_MulAddRecFN.scala 164:35]
  assign mulAddRecFN_io_detectTininess = io_detectTininess; // @[ValExec_MulAddRecFN.scala 165:35]
endmodule
