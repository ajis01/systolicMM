module CompareRecFN(
  input  [32:0] io_a,
  input  [32:0] io_b,
  output        io_lt,
  output        io_eq,
  output [4:0]  io_exceptionFlags
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] rawB_sig; // @[Cat.scala 29:58]
  wire  ordered; // @[CompareRecFN.scala 57:32]
  wire  bothInfs; // @[CompareRecFN.scala 58:33]
  wire  bothZeros; // @[CompareRecFN.scala 59:33]
  wire  eqExps; // @[CompareRecFN.scala 60:29]
  wire  _T_34; // @[CompareRecFN.scala 62:20]
  wire  _T_35; // @[CompareRecFN.scala 62:57]
  wire  _T_36; // @[CompareRecFN.scala 62:44]
  wire  common_ltMags; // @[CompareRecFN.scala 62:33]
  wire  _T_37; // @[CompareRecFN.scala 63:45]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32]
  wire  _T_40; // @[CompareRecFN.scala 67:25]
  wire  _T_43; // @[CompareRecFN.scala 69:35]
  wire  _T_45; // @[CompareRecFN.scala 69:54]
  wire  _T_47; // @[CompareRecFN.scala 70:41]
  wire  _T_48; // @[CompareRecFN.scala 69:74]
  wire  _T_49; // @[CompareRecFN.scala 68:30]
  wire  _T_50; // @[CompareRecFN.scala 67:41]
  wire  ordered_lt; // @[CompareRecFN.scala 66:21]
  wire  _T_51; // @[CompareRecFN.scala 72:34]
  wire  _T_52; // @[CompareRecFN.scala 72:62]
  wire  _T_53; // @[CompareRecFN.scala 72:49]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19]
  wire  _T_56; // @[common.scala 81:46]
  wire  _T_59; // @[common.scala 81:46]
  wire  _T_60; // @[CompareRecFN.scala 75:32]
  wire  invalid; // @[CompareRecFN.scala 75:58]
  assign rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_isInf = _T_4 & ~io_a[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[22:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_isInf = _T_20 & ~io_b[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[22:0]}; // @[Cat.scala 29:58]
  assign ordered = ~rawA_isNaN & ~rawB_isNaN; // @[CompareRecFN.scala 57:32]
  assign bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29]
  assign _T_34 = $signed(rawA_sExp) < $signed(rawB_sExp); // @[CompareRecFN.scala 62:20]
  assign _T_35 = rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:57]
  assign _T_36 = eqExps & _T_35; // @[CompareRecFN.scala 62:44]
  assign common_ltMags = _T_34 | _T_36; // @[CompareRecFN.scala 62:33]
  assign _T_37 = rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:45]
  assign common_eqMags = eqExps & _T_37; // @[CompareRecFN.scala 63:32]
  assign _T_40 = rawA_sign & ~rawB_sign; // @[CompareRecFN.scala 67:25]
  assign _T_43 = rawA_sign & ~common_ltMags; // @[CompareRecFN.scala 69:35]
  assign _T_45 = _T_43 & ~common_eqMags; // @[CompareRecFN.scala 69:54]
  assign _T_47 = ~rawB_sign & common_ltMags; // @[CompareRecFN.scala 70:41]
  assign _T_48 = _T_45 | _T_47; // @[CompareRecFN.scala 69:74]
  assign _T_49 = ~bothInfs & _T_48; // @[CompareRecFN.scala 68:30]
  assign _T_50 = _T_40 | _T_49; // @[CompareRecFN.scala 67:41]
  assign ordered_lt = ~bothZeros & _T_50; // @[CompareRecFN.scala 66:21]
  assign _T_51 = rawA_sign == rawB_sign; // @[CompareRecFN.scala 72:34]
  assign _T_52 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62]
  assign _T_53 = _T_51 & _T_52; // @[CompareRecFN.scala 72:49]
  assign ordered_eq = bothZeros | _T_53; // @[CompareRecFN.scala 72:19]
  assign _T_56 = rawA_isNaN & ~rawA_sig[22]; // @[common.scala 81:46]
  assign _T_59 = rawB_isNaN & ~rawB_sig[22]; // @[common.scala 81:46]
  assign _T_60 = _T_56 | _T_59; // @[CompareRecFN.scala 75:32]
  assign invalid = _T_60 | ~ordered; // @[CompareRecFN.scala 75:58]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:11]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23]
endmodule
module ValExec_CompareRecF32_le(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  input  [31:0] io_b,
  input         io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output        io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [32:0] compareRecFN_io_a; // @[ValExec_CompareRecFN.scala 94:30]
  wire [32:0] compareRecFN_io_b; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 94:30]
  wire [4:0] compareRecFN_io_exceptionFlags; // @[ValExec_CompareRecFN.scala 94:30]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_48; // @[Mux.scala 47:69]
  wire [4:0] _T_49; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61; // @[rawFloatFromFN.scala 63:62]
  wire  _T_64; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_67; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_69; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_71; // @[Cat.scala 29:58]
  wire [2:0] _T_73; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_75; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_78; // @[Cat.scala 29:58]
  wire [3:0] _T_79; // @[Cat.scala 29:58]
  wire  _T_84; // @[rawFloatFromFN.scala 50:34]
  wire  _T_85; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_118; // @[Mux.scala 47:69]
  wire [4:0] _T_119; // @[Mux.scala 47:69]
  wire [4:0] _T_120; // @[Mux.scala 47:69]
  wire [4:0] _T_121; // @[Mux.scala 47:69]
  wire [4:0] _T_122; // @[Mux.scala 47:69]
  wire [4:0] _T_123; // @[Mux.scala 47:69]
  wire [4:0] _T_124; // @[Mux.scala 47:69]
  wire [4:0] _T_125; // @[Mux.scala 47:69]
  wire [4:0] _T_126; // @[Mux.scala 47:69]
  wire [4:0] _T_127; // @[Mux.scala 47:69]
  wire [4:0] _T_128; // @[Mux.scala 47:69]
  wire [4:0] _T_129; // @[Mux.scala 47:69]
  wire [4:0] _T_130; // @[Mux.scala 47:69]
  wire [53:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_131; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_133; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_134; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_135; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_136; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_137; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_139; // @[rawFloatFromFN.scala 59:15]
  wire  _T_140; // @[rawFloatFromFN.scala 62:34]
  wire  _T_142; // @[rawFloatFromFN.scala 63:62]
  wire  _T_145; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_148; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_150; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_152; // @[Cat.scala 29:58]
  wire [2:0] _T_154; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_156; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_159; // @[Cat.scala 29:58]
  wire [3:0] _T_160; // @[Cat.scala 29:58]
  wire  _T_163; // @[ValExec_CompareRecFN.scala 104:24]
  wire  _T_164; // @[ValExec_CompareRecFN.scala 105:35]
  CompareRecFN compareRecFN ( // @[ValExec_CompareRecFN.scala 94:30]
    .io_a(compareRecFN_io_a),
    .io_b(compareRecFN_io_b),
    .io_lt(compareRecFN_io_lt),
    .io_eq(compareRecFN_io_eq),
    .io_exceptionFlags(compareRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  assign _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  assign _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  assign _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  assign _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  assign _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  assign _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  assign _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  assign _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  assign _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  assign _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  assign _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  assign _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  assign _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  assign _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  assign _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  assign _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  assign _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  assign _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  assign _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  assign _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  assign _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  assign _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  assign _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  assign _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  assign _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_64 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_67 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_69 = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_71 = {1'h0,~_T_59,_T_69}; // @[Cat.scala 29:58]
  assign _T_73 = _T_59 ? 3'h0 : _T_67[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_64}; // @[recFNFromFN.scala 48:79]
  assign _T_75 = _T_73 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_78 = {_T_67[5:0],_T_71[22:0]}; // @[Cat.scala 29:58]
  assign _T_79 = {io_a[31],_T_75}; // @[Cat.scala 29:58]
  assign _T_84 = io_b[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_85 = io_b[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_109 = io_b[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_110 = io_b[2] ? 5'h14 : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = io_b[3] ? 5'h13 : _T_110; // @[Mux.scala 47:69]
  assign _T_112 = io_b[4] ? 5'h12 : _T_111; // @[Mux.scala 47:69]
  assign _T_113 = io_b[5] ? 5'h11 : _T_112; // @[Mux.scala 47:69]
  assign _T_114 = io_b[6] ? 5'h10 : _T_113; // @[Mux.scala 47:69]
  assign _T_115 = io_b[7] ? 5'hf : _T_114; // @[Mux.scala 47:69]
  assign _T_116 = io_b[8] ? 5'he : _T_115; // @[Mux.scala 47:69]
  assign _T_117 = io_b[9] ? 5'hd : _T_116; // @[Mux.scala 47:69]
  assign _T_118 = io_b[10] ? 5'hc : _T_117; // @[Mux.scala 47:69]
  assign _T_119 = io_b[11] ? 5'hb : _T_118; // @[Mux.scala 47:69]
  assign _T_120 = io_b[12] ? 5'ha : _T_119; // @[Mux.scala 47:69]
  assign _T_121 = io_b[13] ? 5'h9 : _T_120; // @[Mux.scala 47:69]
  assign _T_122 = io_b[14] ? 5'h8 : _T_121; // @[Mux.scala 47:69]
  assign _T_123 = io_b[15] ? 5'h7 : _T_122; // @[Mux.scala 47:69]
  assign _T_124 = io_b[16] ? 5'h6 : _T_123; // @[Mux.scala 47:69]
  assign _T_125 = io_b[17] ? 5'h5 : _T_124; // @[Mux.scala 47:69]
  assign _T_126 = io_b[18] ? 5'h4 : _T_125; // @[Mux.scala 47:69]
  assign _T_127 = io_b[19] ? 5'h3 : _T_126; // @[Mux.scala 47:69]
  assign _T_128 = io_b[20] ? 5'h2 : _T_127; // @[Mux.scala 47:69]
  assign _T_129 = io_b[21] ? 5'h1 : _T_128; // @[Mux.scala 47:69]
  assign _T_130 = io_b[22] ? 5'h0 : _T_129; // @[Mux.scala 47:69]
  assign _GEN_5 = {{31'd0}, io_b[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_131 = _GEN_5 << _T_130; // @[rawFloatFromFN.scala 54:36]
  assign _T_133 = {_T_131[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{4'd0}, _T_130}; // @[rawFloatFromFN.scala 57:26]
  assign _T_134 = _GEN_6 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_135 = _T_84 ? _T_134 : {{1'd0}, io_b[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_136 = _T_84 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{6'd0}, _T_136}; // @[rawFloatFromFN.scala 60:22]
  assign _T_137 = 8'h80 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_137}; // @[rawFloatFromFN.scala 59:15]
  assign _T_139 = _T_135 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_140 = _T_84 & _T_85; // @[rawFloatFromFN.scala 62:34]
  assign _T_142 = _T_139[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_145 = _T_142 & ~_T_85; // @[rawFloatFromFN.scala 66:33]
  assign _T_148 = {1'b0,$signed(_T_139)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_150 = _T_84 ? _T_133 : io_b[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_152 = {1'h0,~_T_140,_T_150}; // @[Cat.scala 29:58]
  assign _T_154 = _T_140 ? 3'h0 : _T_148[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_145}; // @[recFNFromFN.scala 48:79]
  assign _T_156 = _T_154 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_159 = {_T_148[5:0],_T_152[22:0]}; // @[Cat.scala 29:58]
  assign _T_160 = {io_b[31],_T_156}; // @[Cat.scala 29:58]
  assign _T_163 = io_actual_out == io_expected_out; // @[ValExec_CompareRecFN.scala 104:24]
  assign _T_164 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_CompareRecFN.scala 105:35]
  assign io_actual_out = compareRecFN_io_lt | compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 99:19]
  assign io_actual_exceptionFlags = compareRecFN_io_exceptionFlags; // @[ValExec_CompareRecFN.scala 100:30]
  assign io_check = 1'h1; // @[ValExec_CompareRecFN.scala 102:14]
  assign io_pass = _T_163 & _T_164; // @[ValExec_CompareRecFN.scala 103:13]
  assign compareRecFN_io_a = {_T_79,_T_78}; // @[ValExec_CompareRecFN.scala 95:23]
  assign compareRecFN_io_b = {_T_160,_T_159}; // @[ValExec_CompareRecFN.scala 96:23]
endmodule
