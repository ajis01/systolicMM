module CompareRecFN(
  input  [16:0] io_a,
  input  [16:0] io_b,
  output        io_eq,
  output [4:0]  io_exceptionFlags
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [11:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [11:0] rawB_sig; // @[Cat.scala 29:58]
  wire  ordered; // @[CompareRecFN.scala 57:32]
  wire  bothInfs; // @[CompareRecFN.scala 58:33]
  wire  bothZeros; // @[CompareRecFN.scala 59:33]
  wire  eqExps; // @[CompareRecFN.scala 60:29]
  wire  _T_37; // @[CompareRecFN.scala 63:45]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32]
  wire  _T_51; // @[CompareRecFN.scala 72:34]
  wire  _T_52; // @[CompareRecFN.scala 72:62]
  wire  _T_53; // @[CompareRecFN.scala 72:49]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19]
  wire  _T_56; // @[common.scala 81:46]
  wire  _T_59; // @[common.scala 81:46]
  wire  invalid; // @[CompareRecFN.scala 75:32]
  assign rawA_isZero = io_a[15:13] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[15:14] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[13]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_isInf = _T_4 & ~io_a[13]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA_sign = io_a[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[15:10])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[9:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[15:13] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[15:14] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[13]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_isInf = _T_20 & ~io_b[13]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB_sign = io_b[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[15:10])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[9:0]}; // @[Cat.scala 29:58]
  assign ordered = ~rawA_isNaN & ~rawB_isNaN; // @[CompareRecFN.scala 57:32]
  assign bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29]
  assign _T_37 = rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:45]
  assign common_eqMags = eqExps & _T_37; // @[CompareRecFN.scala 63:32]
  assign _T_51 = rawA_sign == rawB_sign; // @[CompareRecFN.scala 72:34]
  assign _T_52 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62]
  assign _T_53 = _T_51 & _T_52; // @[CompareRecFN.scala 72:49]
  assign ordered_eq = bothZeros | _T_53; // @[CompareRecFN.scala 72:19]
  assign _T_56 = rawA_isNaN & ~rawA_sig[9]; // @[common.scala 81:46]
  assign _T_59 = rawB_isNaN & ~rawB_sig[9]; // @[common.scala 81:46]
  assign invalid = _T_56 | _T_59; // @[CompareRecFN.scala 75:32]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23]
endmodule
module ValExec_CompareRecF16_eq(
  input         clock,
  input         reset,
  input  [15:0] io_a,
  input  [15:0] io_b,
  input         io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output        io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [16:0] compareRecFN_io_a; // @[ValExec_CompareRecFN.scala 129:30]
  wire [16:0] compareRecFN_io_b; // @[ValExec_CompareRecFN.scala 129:30]
  wire  compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 129:30]
  wire [4:0] compareRecFN_io_exceptionFlags; // @[ValExec_CompareRecFN.scala 129:30]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_15; // @[Mux.scala 47:69]
  wire [3:0] _T_16; // @[Mux.scala 47:69]
  wire [3:0] _T_17; // @[Mux.scala 47:69]
  wire [3:0] _T_18; // @[Mux.scala 47:69]
  wire [3:0] _T_19; // @[Mux.scala 47:69]
  wire [3:0] _T_20; // @[Mux.scala 47:69]
  wire [3:0] _T_21; // @[Mux.scala 47:69]
  wire [3:0] _T_22; // @[Mux.scala 47:69]
  wire [3:0] _T_23; // @[Mux.scala 47:69]
  wire [24:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_24; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_26; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_27; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_28; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_29; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_30; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_32; // @[rawFloatFromFN.scala 59:15]
  wire  _T_33; // @[rawFloatFromFN.scala 62:34]
  wire  _T_35; // @[rawFloatFromFN.scala 63:62]
  wire  _T_38; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_41; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_43; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_45; // @[Cat.scala 29:58]
  wire [2:0] _T_47; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_49; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_52; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[Cat.scala 29:58]
  wire  _T_58; // @[rawFloatFromFN.scala 50:34]
  wire  _T_59; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_70; // @[Mux.scala 47:69]
  wire [3:0] _T_71; // @[Mux.scala 47:69]
  wire [3:0] _T_72; // @[Mux.scala 47:69]
  wire [3:0] _T_73; // @[Mux.scala 47:69]
  wire [3:0] _T_74; // @[Mux.scala 47:69]
  wire [3:0] _T_75; // @[Mux.scala 47:69]
  wire [3:0] _T_76; // @[Mux.scala 47:69]
  wire [3:0] _T_77; // @[Mux.scala 47:69]
  wire [3:0] _T_78; // @[Mux.scala 47:69]
  wire [24:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_79; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_81; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_82; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_83; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_84; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_85; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_87; // @[rawFloatFromFN.scala 59:15]
  wire  _T_88; // @[rawFloatFromFN.scala 62:34]
  wire  _T_90; // @[rawFloatFromFN.scala 63:62]
  wire  _T_93; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_96; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_98; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_100; // @[Cat.scala 29:58]
  wire [2:0] _T_102; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_104; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_107; // @[Cat.scala 29:58]
  wire [3:0] _T_108; // @[Cat.scala 29:58]
  wire  _T_110; // @[ValExec_CompareRecFN.scala 139:24]
  wire  _T_111; // @[ValExec_CompareRecFN.scala 140:35]
  CompareRecFN compareRecFN ( // @[ValExec_CompareRecFN.scala 129:30]
    .io_a(compareRecFN_io_a),
    .io_b(compareRecFN_io_b),
    .io_eq(compareRecFN_io_eq),
    .io_exceptionFlags(compareRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_a[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_a[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_15 = io_a[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_16 = io_a[2] ? 4'h7 : _T_15; // @[Mux.scala 47:69]
  assign _T_17 = io_a[3] ? 4'h6 : _T_16; // @[Mux.scala 47:69]
  assign _T_18 = io_a[4] ? 4'h5 : _T_17; // @[Mux.scala 47:69]
  assign _T_19 = io_a[5] ? 4'h4 : _T_18; // @[Mux.scala 47:69]
  assign _T_20 = io_a[6] ? 4'h3 : _T_19; // @[Mux.scala 47:69]
  assign _T_21 = io_a[7] ? 4'h2 : _T_20; // @[Mux.scala 47:69]
  assign _T_22 = io_a[8] ? 4'h1 : _T_21; // @[Mux.scala 47:69]
  assign _T_23 = io_a[9] ? 4'h0 : _T_22; // @[Mux.scala 47:69]
  assign _GEN_0 = {{15'd0}, io_a[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_24 = _GEN_0 << _T_23; // @[rawFloatFromFN.scala 54:36]
  assign _T_26 = {_T_24[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{2'd0}, _T_23}; // @[rawFloatFromFN.scala 57:26]
  assign _T_27 = _GEN_1 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_28 = _T_3 ? _T_27 : {{1'd0}, io_a[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_29 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{3'd0}, _T_29}; // @[rawFloatFromFN.scala 60:22]
  assign _T_30 = 5'h10 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_30}; // @[rawFloatFromFN.scala 59:15]
  assign _T_32 = _T_28 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_33 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_35 = _T_32[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_38 = _T_35 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_41 = {1'b0,$signed(_T_32)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_43 = _T_3 ? _T_26 : io_a[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_45 = {1'h0,~_T_33,_T_43}; // @[Cat.scala 29:58]
  assign _T_47 = _T_33 ? 3'h0 : _T_41[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_38}; // @[recFNFromFN.scala 48:79]
  assign _T_49 = _T_47 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_52 = {_T_41[2:0],_T_45[9:0]}; // @[Cat.scala 29:58]
  assign _T_53 = {io_a[15],_T_49}; // @[Cat.scala 29:58]
  assign _T_58 = io_b[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_59 = io_b[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_70 = io_b[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_71 = io_b[2] ? 4'h7 : _T_70; // @[Mux.scala 47:69]
  assign _T_72 = io_b[3] ? 4'h6 : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = io_b[4] ? 4'h5 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = io_b[5] ? 4'h4 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = io_b[6] ? 4'h3 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = io_b[7] ? 4'h2 : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = io_b[8] ? 4'h1 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = io_b[9] ? 4'h0 : _T_77; // @[Mux.scala 47:69]
  assign _GEN_5 = {{15'd0}, io_b[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_79 = _GEN_5 << _T_78; // @[rawFloatFromFN.scala 54:36]
  assign _T_81 = {_T_79[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{2'd0}, _T_78}; // @[rawFloatFromFN.scala 57:26]
  assign _T_82 = _GEN_6 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_83 = _T_58 ? _T_82 : {{1'd0}, io_b[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_84 = _T_58 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{3'd0}, _T_84}; // @[rawFloatFromFN.scala 60:22]
  assign _T_85 = 5'h10 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_85}; // @[rawFloatFromFN.scala 59:15]
  assign _T_87 = _T_83 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_88 = _T_58 & _T_59; // @[rawFloatFromFN.scala 62:34]
  assign _T_90 = _T_87[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_93 = _T_90 & ~_T_59; // @[rawFloatFromFN.scala 66:33]
  assign _T_96 = {1'b0,$signed(_T_87)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_98 = _T_58 ? _T_81 : io_b[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_100 = {1'h0,~_T_88,_T_98}; // @[Cat.scala 29:58]
  assign _T_102 = _T_88 ? 3'h0 : _T_96[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_93}; // @[recFNFromFN.scala 48:79]
  assign _T_104 = _T_102 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_107 = {_T_96[2:0],_T_100[9:0]}; // @[Cat.scala 29:58]
  assign _T_108 = {io_b[15],_T_104}; // @[Cat.scala 29:58]
  assign _T_110 = io_actual_out == io_expected_out; // @[ValExec_CompareRecFN.scala 139:24]
  assign _T_111 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_CompareRecFN.scala 140:35]
  assign io_actual_out = compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 134:19]
  assign io_actual_exceptionFlags = compareRecFN_io_exceptionFlags; // @[ValExec_CompareRecFN.scala 135:30]
  assign io_check = 1'h1; // @[ValExec_CompareRecFN.scala 137:14]
  assign io_pass = _T_110 & _T_111; // @[ValExec_CompareRecFN.scala 138:13]
  assign compareRecFN_io_a = {_T_53,_T_52}; // @[ValExec_CompareRecFN.scala 130:23]
  assign compareRecFN_io_b = {_T_108,_T_107}; // @[ValExec_CompareRecFN.scala 131:23]
endmodule
