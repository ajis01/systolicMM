module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [24:0] io_in_sig,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire [11:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] _T_3; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire [55:0] adjustedSig; // @[RoundAnyRawFNToRecFN.scala 112:22]
  wire [12:0] _T_6; // @[RoundAnyRawFNToRecFN.scala 134:55]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 134:55]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 138:28]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire [11:0] _T_22; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _T_24; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [11:0] _T_32; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [11:0] _T_34; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [11:0] _T_39; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [11:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [11:0] _T_41; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_42; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire [51:0] _T_44; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [12:0] _T_48; // @[Cat.scala 29:58]
  wire [2:0] _T_52; // @[Cat.scala 29:58]
  assign _GEN_0 = {{2{io_in_sExp[9]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign _T_3 = $signed(_GEN_0) + 12'sh700; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_T_3[11:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign adjustedSig = {io_in_sig, 31'h0}; // @[RoundAnyRawFNToRecFN.scala 112:22]
  assign _T_6 = {{1'd0}, sAdjustedExp[11:0]}; // @[RoundAnyRawFNToRecFN.scala 134:55]
  assign common_expOut = _T_6[11:0]; // @[RoundAnyRawFNToRecFN.scala 134:55]
  assign common_fractOut = adjustedSig[53:2]; // @[RoundAnyRawFNToRecFN.scala 138:28]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_22 = io_in_isZero ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_24 = common_expOut & ~_T_22; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_32 = io_in_isInf ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_34 = _T_24 & ~_T_32; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_39 = io_in_isInf ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_40 = _T_34 | _T_39; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_41 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_40 | _T_41; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_42 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_44 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign fractOut = _T_42 ? _T_44 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_48 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_52 = {io_invalidExc,1'h0,1'h0}; // @[Cat.scala 29:58]
  assign io_out = {_T_48,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_52,2'h0}; // @[RoundAnyRawFNToRecFN.scala 285:23]
endmodule
module RecFNToRecFN(
  input  [32:0] io_in,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  RoundAnyRawFNToRecFN_io_invalidExc; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isNaN; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isInf; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isZero; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_sign; // @[RecFNToRecFN.scala 72:19]
  wire [9:0] RoundAnyRawFNToRecFN_io_in_sExp; // @[RecFNToRecFN.scala 72:19]
  wire [24:0] RoundAnyRawFNToRecFN_io_in_sig; // @[RecFNToRecFN.scala 72:19]
  wire [64:0] RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 72:19]
  wire [4:0] RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 72:19]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [24:0] rawIn_sig; // @[Cat.scala 29:58]
  RoundAnyRawFNToRecFN RoundAnyRawFNToRecFN ( // @[RecFNToRecFN.scala 72:19]
    .io_invalidExc(RoundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(RoundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(RoundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(RoundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(RoundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(RoundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(RoundAnyRawFNToRecFN_io_in_sig),
    .io_out(RoundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(RoundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign rawIn_isZero = io_in[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_in[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_4 & io_in[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_14 = {1'h0,~rawIn_isZero}; // @[Cat.scala 29:58]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[22:0]}; // @[Cat.scala 29:58]
  assign io_out = RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 85:27]
  assign io_exceptionFlags = RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 86:27]
  assign RoundAnyRawFNToRecFN_io_invalidExc = rawIn_isNaN & ~rawIn_sig[22]; // @[RecFNToRecFN.scala 80:48]
  assign RoundAnyRawFNToRecFN_io_in_isNaN = _T_4 & io_in[29]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isInf = _T_4 & ~io_in[29]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isZero = io_in[31:29] == 3'h0; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sign = io_in[32]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(io_in[31:23])}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sig = {_T_14,io_in[22:0]}; // @[RecFNToRecFN.scala 82:48]
endmodule
module ValExec_RecF32ToRecF64(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [63:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [64:0] io_expected_recOut,
  output [64:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [32:0] recFNToRecFN_io_in; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire [64:0] recFNToRecFN_io_out; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire [4:0] recFNToRecFN_io_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_48; // @[Mux.scala 47:69]
  wire [4:0] _T_49; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61; // @[rawFloatFromFN.scala 63:62]
  wire  _T_64; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_67; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_69; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_71; // @[Cat.scala 29:58]
  wire [2:0] _T_73; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_75; // @[recFNFromFN.scala 48:79]
  wire [28:0] _T_78; // @[Cat.scala 29:58]
  wire [3:0] _T_79; // @[Cat.scala 29:58]
  wire  _T_84; // @[rawFloatFromFN.scala 50:34]
  wire  _T_85; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_138; // @[Mux.scala 47:69]
  wire [5:0] _T_139; // @[Mux.scala 47:69]
  wire [5:0] _T_140; // @[Mux.scala 47:69]
  wire [5:0] _T_141; // @[Mux.scala 47:69]
  wire [5:0] _T_142; // @[Mux.scala 47:69]
  wire [5:0] _T_143; // @[Mux.scala 47:69]
  wire [5:0] _T_144; // @[Mux.scala 47:69]
  wire [5:0] _T_145; // @[Mux.scala 47:69]
  wire [5:0] _T_146; // @[Mux.scala 47:69]
  wire [5:0] _T_147; // @[Mux.scala 47:69]
  wire [5:0] _T_148; // @[Mux.scala 47:69]
  wire [5:0] _T_149; // @[Mux.scala 47:69]
  wire [5:0] _T_150; // @[Mux.scala 47:69]
  wire [5:0] _T_151; // @[Mux.scala 47:69]
  wire [5:0] _T_152; // @[Mux.scala 47:69]
  wire [5:0] _T_153; // @[Mux.scala 47:69]
  wire [5:0] _T_154; // @[Mux.scala 47:69]
  wire [5:0] _T_155; // @[Mux.scala 47:69]
  wire [5:0] _T_156; // @[Mux.scala 47:69]
  wire [5:0] _T_157; // @[Mux.scala 47:69]
  wire [5:0] _T_158; // @[Mux.scala 47:69]
  wire [5:0] _T_159; // @[Mux.scala 47:69]
  wire [5:0] _T_160; // @[Mux.scala 47:69]
  wire [5:0] _T_161; // @[Mux.scala 47:69]
  wire [5:0] _T_162; // @[Mux.scala 47:69]
  wire [5:0] _T_163; // @[Mux.scala 47:69]
  wire [5:0] _T_164; // @[Mux.scala 47:69]
  wire [5:0] _T_165; // @[Mux.scala 47:69]
  wire [5:0] _T_166; // @[Mux.scala 47:69]
  wire [5:0] _T_167; // @[Mux.scala 47:69]
  wire [5:0] _T_168; // @[Mux.scala 47:69]
  wire [5:0] _T_169; // @[Mux.scala 47:69]
  wire [5:0] _T_170; // @[Mux.scala 47:69]
  wire [5:0] _T_171; // @[Mux.scala 47:69]
  wire [5:0] _T_172; // @[Mux.scala 47:69]
  wire [5:0] _T_173; // @[Mux.scala 47:69]
  wire [5:0] _T_174; // @[Mux.scala 47:69]
  wire [5:0] _T_175; // @[Mux.scala 47:69]
  wire [5:0] _T_176; // @[Mux.scala 47:69]
  wire [5:0] _T_177; // @[Mux.scala 47:69]
  wire [5:0] _T_178; // @[Mux.scala 47:69]
  wire [5:0] _T_179; // @[Mux.scala 47:69]
  wire [5:0] _T_180; // @[Mux.scala 47:69]
  wire [5:0] _T_181; // @[Mux.scala 47:69]
  wire [5:0] _T_182; // @[Mux.scala 47:69]
  wire [5:0] _T_183; // @[Mux.scala 47:69]
  wire [5:0] _T_184; // @[Mux.scala 47:69]
  wire [5:0] _T_185; // @[Mux.scala 47:69]
  wire [5:0] _T_186; // @[Mux.scala 47:69]
  wire [5:0] _T_187; // @[Mux.scala 47:69]
  wire [5:0] _T_188; // @[Mux.scala 47:69]
  wire [114:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_189; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_191; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_192; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_193; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_194; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_195; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_197; // @[rawFloatFromFN.scala 59:15]
  wire  _T_198; // @[rawFloatFromFN.scala 62:34]
  wire  _T_200; // @[rawFloatFromFN.scala 63:62]
  wire  _T_203; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_206; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_208; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_210; // @[Cat.scala 29:58]
  wire [2:0] _T_212; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_214; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_217; // @[Cat.scala 29:58]
  wire [3:0] _T_218; // @[Cat.scala 29:58]
  wire  _T_223; // @[tests.scala 48:26]
  wire  _T_225; // @[tests.scala 48:55]
  wire  _T_226; // @[tests.scala 48:39]
  wire  _T_227; // @[tests.scala 49:20]
  wire  _T_230; // @[tests.scala 49:54]
  wire  _T_231; // @[tests.scala 49:31]
  wire  _T_233; // @[tests.scala 50:30]
  wire  _T_235; // @[tests.scala 50:66]
  wire  _T_236; // @[tests.scala 50:16]
  wire  _T_237; // @[tests.scala 48:12]
  wire  _T_238; // @[ValExec_RecFNToRecFN.scala 84:35]
  RecFNToRecFN recFNToRecFN ( // @[ValExec_RecFNToRecFN.scala 68:15]
    .io_in(recFNToRecFN_io_in),
    .io_out(recFNToRecFN_io_out),
    .io_exceptionFlags(recFNToRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_in[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_in[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_28 = io_in[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_29 = io_in[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  assign _T_30 = io_in[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  assign _T_31 = io_in[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  assign _T_32 = io_in[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  assign _T_33 = io_in[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  assign _T_34 = io_in[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  assign _T_35 = io_in[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  assign _T_36 = io_in[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  assign _T_37 = io_in[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  assign _T_38 = io_in[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  assign _T_39 = io_in[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  assign _T_40 = io_in[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  assign _T_41 = io_in[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  assign _T_42 = io_in[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  assign _T_43 = io_in[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  assign _T_44 = io_in[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  assign _T_45 = io_in[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  assign _T_46 = io_in[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  assign _T_47 = io_in[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  assign _T_48 = io_in[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  assign _T_49 = io_in[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  assign _GEN_0 = {{31'd0}, io_in[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  assign _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  assign _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_54 = _T_3 ? _T_53 : {{1'd0}, io_in[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  assign _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  assign _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_64 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_67 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_69 = _T_3 ? _T_52 : io_in[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_71 = {1'h0,~_T_59,_T_69}; // @[Cat.scala 29:58]
  assign _T_73 = _T_59 ? 3'h0 : _T_67[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_64}; // @[recFNFromFN.scala 48:79]
  assign _T_75 = _T_73 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_78 = {_T_67[5:0],_T_71[22:0]}; // @[Cat.scala 29:58]
  assign _T_79 = {io_in[31],_T_75}; // @[Cat.scala 29:58]
  assign _T_84 = io_expected_out[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_85 = io_expected_out[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_138 = io_expected_out[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_139 = io_expected_out[2] ? 6'h31 : _T_138; // @[Mux.scala 47:69]
  assign _T_140 = io_expected_out[3] ? 6'h30 : _T_139; // @[Mux.scala 47:69]
  assign _T_141 = io_expected_out[4] ? 6'h2f : _T_140; // @[Mux.scala 47:69]
  assign _T_142 = io_expected_out[5] ? 6'h2e : _T_141; // @[Mux.scala 47:69]
  assign _T_143 = io_expected_out[6] ? 6'h2d : _T_142; // @[Mux.scala 47:69]
  assign _T_144 = io_expected_out[7] ? 6'h2c : _T_143; // @[Mux.scala 47:69]
  assign _T_145 = io_expected_out[8] ? 6'h2b : _T_144; // @[Mux.scala 47:69]
  assign _T_146 = io_expected_out[9] ? 6'h2a : _T_145; // @[Mux.scala 47:69]
  assign _T_147 = io_expected_out[10] ? 6'h29 : _T_146; // @[Mux.scala 47:69]
  assign _T_148 = io_expected_out[11] ? 6'h28 : _T_147; // @[Mux.scala 47:69]
  assign _T_149 = io_expected_out[12] ? 6'h27 : _T_148; // @[Mux.scala 47:69]
  assign _T_150 = io_expected_out[13] ? 6'h26 : _T_149; // @[Mux.scala 47:69]
  assign _T_151 = io_expected_out[14] ? 6'h25 : _T_150; // @[Mux.scala 47:69]
  assign _T_152 = io_expected_out[15] ? 6'h24 : _T_151; // @[Mux.scala 47:69]
  assign _T_153 = io_expected_out[16] ? 6'h23 : _T_152; // @[Mux.scala 47:69]
  assign _T_154 = io_expected_out[17] ? 6'h22 : _T_153; // @[Mux.scala 47:69]
  assign _T_155 = io_expected_out[18] ? 6'h21 : _T_154; // @[Mux.scala 47:69]
  assign _T_156 = io_expected_out[19] ? 6'h20 : _T_155; // @[Mux.scala 47:69]
  assign _T_157 = io_expected_out[20] ? 6'h1f : _T_156; // @[Mux.scala 47:69]
  assign _T_158 = io_expected_out[21] ? 6'h1e : _T_157; // @[Mux.scala 47:69]
  assign _T_159 = io_expected_out[22] ? 6'h1d : _T_158; // @[Mux.scala 47:69]
  assign _T_160 = io_expected_out[23] ? 6'h1c : _T_159; // @[Mux.scala 47:69]
  assign _T_161 = io_expected_out[24] ? 6'h1b : _T_160; // @[Mux.scala 47:69]
  assign _T_162 = io_expected_out[25] ? 6'h1a : _T_161; // @[Mux.scala 47:69]
  assign _T_163 = io_expected_out[26] ? 6'h19 : _T_162; // @[Mux.scala 47:69]
  assign _T_164 = io_expected_out[27] ? 6'h18 : _T_163; // @[Mux.scala 47:69]
  assign _T_165 = io_expected_out[28] ? 6'h17 : _T_164; // @[Mux.scala 47:69]
  assign _T_166 = io_expected_out[29] ? 6'h16 : _T_165; // @[Mux.scala 47:69]
  assign _T_167 = io_expected_out[30] ? 6'h15 : _T_166; // @[Mux.scala 47:69]
  assign _T_168 = io_expected_out[31] ? 6'h14 : _T_167; // @[Mux.scala 47:69]
  assign _T_169 = io_expected_out[32] ? 6'h13 : _T_168; // @[Mux.scala 47:69]
  assign _T_170 = io_expected_out[33] ? 6'h12 : _T_169; // @[Mux.scala 47:69]
  assign _T_171 = io_expected_out[34] ? 6'h11 : _T_170; // @[Mux.scala 47:69]
  assign _T_172 = io_expected_out[35] ? 6'h10 : _T_171; // @[Mux.scala 47:69]
  assign _T_173 = io_expected_out[36] ? 6'hf : _T_172; // @[Mux.scala 47:69]
  assign _T_174 = io_expected_out[37] ? 6'he : _T_173; // @[Mux.scala 47:69]
  assign _T_175 = io_expected_out[38] ? 6'hd : _T_174; // @[Mux.scala 47:69]
  assign _T_176 = io_expected_out[39] ? 6'hc : _T_175; // @[Mux.scala 47:69]
  assign _T_177 = io_expected_out[40] ? 6'hb : _T_176; // @[Mux.scala 47:69]
  assign _T_178 = io_expected_out[41] ? 6'ha : _T_177; // @[Mux.scala 47:69]
  assign _T_179 = io_expected_out[42] ? 6'h9 : _T_178; // @[Mux.scala 47:69]
  assign _T_180 = io_expected_out[43] ? 6'h8 : _T_179; // @[Mux.scala 47:69]
  assign _T_181 = io_expected_out[44] ? 6'h7 : _T_180; // @[Mux.scala 47:69]
  assign _T_182 = io_expected_out[45] ? 6'h6 : _T_181; // @[Mux.scala 47:69]
  assign _T_183 = io_expected_out[46] ? 6'h5 : _T_182; // @[Mux.scala 47:69]
  assign _T_184 = io_expected_out[47] ? 6'h4 : _T_183; // @[Mux.scala 47:69]
  assign _T_185 = io_expected_out[48] ? 6'h3 : _T_184; // @[Mux.scala 47:69]
  assign _T_186 = io_expected_out[49] ? 6'h2 : _T_185; // @[Mux.scala 47:69]
  assign _T_187 = io_expected_out[50] ? 6'h1 : _T_186; // @[Mux.scala 47:69]
  assign _T_188 = io_expected_out[51] ? 6'h0 : _T_187; // @[Mux.scala 47:69]
  assign _GEN_5 = {{63'd0}, io_expected_out[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_189 = _GEN_5 << _T_188; // @[rawFloatFromFN.scala 54:36]
  assign _T_191 = {_T_189[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{6'd0}, _T_188}; // @[rawFloatFromFN.scala 57:26]
  assign _T_192 = _GEN_6 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_193 = _T_84 ? _T_192 : {{1'd0}, io_expected_out[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_194 = _T_84 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{9'd0}, _T_194}; // @[rawFloatFromFN.scala 60:22]
  assign _T_195 = 11'h400 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_195}; // @[rawFloatFromFN.scala 59:15]
  assign _T_197 = _T_193 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_198 = _T_84 & _T_85; // @[rawFloatFromFN.scala 62:34]
  assign _T_200 = _T_197[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_203 = _T_200 & ~_T_85; // @[rawFloatFromFN.scala 66:33]
  assign _T_206 = {1'b0,$signed(_T_197)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_208 = _T_84 ? _T_191 : io_expected_out[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_210 = {1'h0,~_T_198,_T_208}; // @[Cat.scala 29:58]
  assign _T_212 = _T_198 ? 3'h0 : _T_206[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_203}; // @[recFNFromFN.scala 48:79]
  assign _T_214 = _T_212 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_217 = {_T_206[8:0],_T_210[51:0]}; // @[Cat.scala 29:58]
  assign _T_218 = {io_expected_out[63],_T_214}; // @[Cat.scala 29:58]
  assign _T_223 = io_actual_out[63:61] == 3'h0; // @[tests.scala 48:26]
  assign _T_225 = io_actual_out[63:61] == 3'h7; // @[tests.scala 48:55]
  assign _T_226 = _T_223 | _T_225; // @[tests.scala 48:39]
  assign _T_227 = io_actual_out[64:61] == io_expected_recOut[64:61]; // @[tests.scala 49:20]
  assign _T_230 = io_actual_out[51:0] == io_expected_recOut[51:0]; // @[tests.scala 49:54]
  assign _T_231 = _T_227 & _T_230; // @[tests.scala 49:31]
  assign _T_233 = io_actual_out[63:61] == 3'h6; // @[tests.scala 50:30]
  assign _T_235 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_236 = _T_233 ? _T_227 : _T_235; // @[tests.scala 50:16]
  assign _T_237 = _T_226 ? _T_231 : _T_236; // @[tests.scala 48:12]
  assign _T_238 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 84:35]
  assign io_expected_recOut = {_T_218,_T_217}; // @[ValExec_RecFNToRecFN.scala 74:24]
  assign io_actual_out = recFNToRecFN_io_out; // @[ValExec_RecFNToRecFN.scala 77:19]
  assign io_actual_exceptionFlags = recFNToRecFN_io_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 78:30]
  assign io_check = 1'h1; // @[ValExec_RecFNToRecFN.scala 80:14]
  assign io_pass = _T_237 & _T_238; // @[ValExec_RecFNToRecFN.scala 81:13]
  assign recFNToRecFN_io_in = {_T_79,_T_78}; // @[ValExec_RecFNToRecFN.scala 70:24]
endmodule
