module ValExec_f32FromRecF32(
  input         clock,
  input         reset,
  input  [31:0] io_a,
  output [31:0] io_out,
  output        io_check,
  output        io_pass
);
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _T_28; // @[Mux.scala 47:69]
  wire [4:0] _T_29; // @[Mux.scala 47:69]
  wire [4:0] _T_30; // @[Mux.scala 47:69]
  wire [4:0] _T_31; // @[Mux.scala 47:69]
  wire [4:0] _T_32; // @[Mux.scala 47:69]
  wire [4:0] _T_33; // @[Mux.scala 47:69]
  wire [4:0] _T_34; // @[Mux.scala 47:69]
  wire [4:0] _T_35; // @[Mux.scala 47:69]
  wire [4:0] _T_36; // @[Mux.scala 47:69]
  wire [4:0] _T_37; // @[Mux.scala 47:69]
  wire [4:0] _T_38; // @[Mux.scala 47:69]
  wire [4:0] _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_48; // @[Mux.scala 47:69]
  wire [4:0] _T_49; // @[Mux.scala 47:69]
  wire [53:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _T_50; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] _T_52; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_53; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _T_54; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_55; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _T_56; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] _T_58; // @[rawFloatFromFN.scala 59:15]
  wire  _T_59; // @[rawFloatFromFN.scala 62:34]
  wire  _T_61; // @[rawFloatFromFN.scala 63:62]
  wire  _T_64; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] _T_67; // @[rawFloatFromFN.scala 70:48]
  wire [22:0] _T_69; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] _T_71; // @[Cat.scala 29:58]
  wire [2:0] _T_73; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_75; // @[recFNFromFN.scala 48:79]
  wire [32:0] _T_80; // @[Cat.scala 29:58]
  wire  _T_83; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_85; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_88; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_91; // @[rawFloatFromRecFN.scala 56:33]
  wire [9:0] _T_93; // @[rawFloatFromRecFN.scala 59:27]
  wire [24:0] _T_97; // @[Cat.scala 29:58]
  wire  _T_98; // @[fNFromRecFN.scala 50:39]
  wire [4:0] _T_101; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _T_103; // @[fNFromRecFN.scala 52:42]
  wire [7:0] _T_107; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _T_108; // @[fNFromRecFN.scala 55:16]
  wire  _T_109; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _T_111; // @[Bitwise.scala 71:12]
  wire [7:0] _T_112; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _T_114; // @[fNFromRecFN.scala 63:20]
  wire [22:0] _T_115; // @[fNFromRecFN.scala 61:16]
  wire [8:0] _T_116; // @[Cat.scala 29:58]
  assign _T_3 = io_a[30:23] == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_a[22:0] == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_28 = io_a[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _T_29 = io_a[2] ? 5'h14 : _T_28; // @[Mux.scala 47:69]
  assign _T_30 = io_a[3] ? 5'h13 : _T_29; // @[Mux.scala 47:69]
  assign _T_31 = io_a[4] ? 5'h12 : _T_30; // @[Mux.scala 47:69]
  assign _T_32 = io_a[5] ? 5'h11 : _T_31; // @[Mux.scala 47:69]
  assign _T_33 = io_a[6] ? 5'h10 : _T_32; // @[Mux.scala 47:69]
  assign _T_34 = io_a[7] ? 5'hf : _T_33; // @[Mux.scala 47:69]
  assign _T_35 = io_a[8] ? 5'he : _T_34; // @[Mux.scala 47:69]
  assign _T_36 = io_a[9] ? 5'hd : _T_35; // @[Mux.scala 47:69]
  assign _T_37 = io_a[10] ? 5'hc : _T_36; // @[Mux.scala 47:69]
  assign _T_38 = io_a[11] ? 5'hb : _T_37; // @[Mux.scala 47:69]
  assign _T_39 = io_a[12] ? 5'ha : _T_38; // @[Mux.scala 47:69]
  assign _T_40 = io_a[13] ? 5'h9 : _T_39; // @[Mux.scala 47:69]
  assign _T_41 = io_a[14] ? 5'h8 : _T_40; // @[Mux.scala 47:69]
  assign _T_42 = io_a[15] ? 5'h7 : _T_41; // @[Mux.scala 47:69]
  assign _T_43 = io_a[16] ? 5'h6 : _T_42; // @[Mux.scala 47:69]
  assign _T_44 = io_a[17] ? 5'h5 : _T_43; // @[Mux.scala 47:69]
  assign _T_45 = io_a[18] ? 5'h4 : _T_44; // @[Mux.scala 47:69]
  assign _T_46 = io_a[19] ? 5'h3 : _T_45; // @[Mux.scala 47:69]
  assign _T_47 = io_a[20] ? 5'h2 : _T_46; // @[Mux.scala 47:69]
  assign _T_48 = io_a[21] ? 5'h1 : _T_47; // @[Mux.scala 47:69]
  assign _T_49 = io_a[22] ? 5'h0 : _T_48; // @[Mux.scala 47:69]
  assign _GEN_0 = {{31'd0}, io_a[22:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_50 = _GEN_0 << _T_49; // @[rawFloatFromFN.scala 54:36]
  assign _T_52 = {_T_50[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{4'd0}, _T_49}; // @[rawFloatFromFN.scala 57:26]
  assign _T_53 = _GEN_1 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _T_54 = _T_3 ? _T_53 : {{1'd0}, io_a[30:23]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_55 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{6'd0}, _T_55}; // @[rawFloatFromFN.scala 60:22]
  assign _T_56 = 8'h80 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_56}; // @[rawFloatFromFN.scala 59:15]
  assign _T_58 = _T_54 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_59 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_61 = _T_58[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_64 = _T_61 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_67 = {1'b0,$signed(_T_58)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_69 = _T_3 ? _T_52 : io_a[22:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_71 = {1'h0,~_T_59,_T_69}; // @[Cat.scala 29:58]
  assign _T_73 = _T_59 ? 3'h0 : _T_67[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_64}; // @[recFNFromFN.scala 48:79]
  assign _T_75 = _T_73 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_80 = {io_a[31],_T_75,_T_67[5:0],_T_71[22:0]}; // @[Cat.scala 29:58]
  assign _T_83 = _T_80[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_85 = _T_80[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign _T_88 = _T_85 & _T_80[29]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_91 = _T_85 & ~_T_80[29]; // @[rawFloatFromRecFN.scala 56:33]
  assign _T_93 = {1'b0,$signed(_T_80[31:23])}; // @[rawFloatFromRecFN.scala 59:27]
  assign _T_97 = {1'h0,~_T_83,_T_80[22:0]}; // @[Cat.scala 29:58]
  assign _T_98 = $signed(_T_93) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  assign _T_101 = 5'h1 - _T_93[4:0]; // @[fNFromRecFN.scala 51:39]
  assign _T_103 = _T_97[24:1] >> _T_101; // @[fNFromRecFN.scala 52:42]
  assign _T_107 = _T_93[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  assign _T_108 = _T_98 ? 8'h0 : _T_107; // @[fNFromRecFN.scala 55:16]
  assign _T_109 = _T_88 | _T_91; // @[fNFromRecFN.scala 59:44]
  assign _T_111 = _T_109 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_112 = _T_108 | _T_111; // @[fNFromRecFN.scala 59:15]
  assign _T_114 = _T_91 ? 23'h0 : _T_97[22:0]; // @[fNFromRecFN.scala 63:20]
  assign _T_115 = _T_98 ? _T_103[22:0] : _T_114; // @[fNFromRecFN.scala 61:16]
  assign _T_116 = {_T_80[32],_T_112}; // @[Cat.scala 29:58]
  assign io_out = {_T_116,_T_115}; // @[ValExec_fNFromRecFN.scala 51:12]
  assign io_check = 1'h1; // @[ValExec_fNFromRecFN.scala 54:14]
  assign io_pass = io_out == io_a; // @[ValExec_fNFromRecFN.scala 55:13]
endmodule
