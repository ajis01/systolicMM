module CompareRecFN(
  input  [64:0] io_a,
  input  [64:0] io_b,
  output        io_lt,
  output        io_eq,
  output [4:0]  io_exceptionFlags
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [53:0] rawB_sig; // @[Cat.scala 29:58]
  wire  ordered; // @[CompareRecFN.scala 57:32]
  wire  bothInfs; // @[CompareRecFN.scala 58:33]
  wire  bothZeros; // @[CompareRecFN.scala 59:33]
  wire  eqExps; // @[CompareRecFN.scala 60:29]
  wire  _T_34; // @[CompareRecFN.scala 62:20]
  wire  _T_35; // @[CompareRecFN.scala 62:57]
  wire  _T_36; // @[CompareRecFN.scala 62:44]
  wire  common_ltMags; // @[CompareRecFN.scala 62:33]
  wire  _T_37; // @[CompareRecFN.scala 63:45]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32]
  wire  _T_40; // @[CompareRecFN.scala 67:25]
  wire  _T_43; // @[CompareRecFN.scala 69:35]
  wire  _T_45; // @[CompareRecFN.scala 69:54]
  wire  _T_47; // @[CompareRecFN.scala 70:41]
  wire  _T_48; // @[CompareRecFN.scala 69:74]
  wire  _T_49; // @[CompareRecFN.scala 68:30]
  wire  _T_50; // @[CompareRecFN.scala 67:41]
  wire  ordered_lt; // @[CompareRecFN.scala 66:21]
  wire  _T_51; // @[CompareRecFN.scala 72:34]
  wire  _T_52; // @[CompareRecFN.scala 72:62]
  wire  _T_53; // @[CompareRecFN.scala 72:49]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19]
  wire  _T_56; // @[common.scala 81:46]
  wire  _T_59; // @[common.scala 81:46]
  wire  _T_60; // @[CompareRecFN.scala 75:32]
  wire  invalid; // @[CompareRecFN.scala 75:58]
  assign rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_isInf = _T_4 & ~io_a[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[51:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_isInf = _T_20 & ~io_b[61]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[51:0]}; // @[Cat.scala 29:58]
  assign ordered = ~rawA_isNaN & ~rawB_isNaN; // @[CompareRecFN.scala 57:32]
  assign bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29]
  assign _T_34 = $signed(rawA_sExp) < $signed(rawB_sExp); // @[CompareRecFN.scala 62:20]
  assign _T_35 = rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:57]
  assign _T_36 = eqExps & _T_35; // @[CompareRecFN.scala 62:44]
  assign common_ltMags = _T_34 | _T_36; // @[CompareRecFN.scala 62:33]
  assign _T_37 = rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:45]
  assign common_eqMags = eqExps & _T_37; // @[CompareRecFN.scala 63:32]
  assign _T_40 = rawA_sign & ~rawB_sign; // @[CompareRecFN.scala 67:25]
  assign _T_43 = rawA_sign & ~common_ltMags; // @[CompareRecFN.scala 69:35]
  assign _T_45 = _T_43 & ~common_eqMags; // @[CompareRecFN.scala 69:54]
  assign _T_47 = ~rawB_sign & common_ltMags; // @[CompareRecFN.scala 70:41]
  assign _T_48 = _T_45 | _T_47; // @[CompareRecFN.scala 69:74]
  assign _T_49 = ~bothInfs & _T_48; // @[CompareRecFN.scala 68:30]
  assign _T_50 = _T_40 | _T_49; // @[CompareRecFN.scala 67:41]
  assign ordered_lt = ~bothZeros & _T_50; // @[CompareRecFN.scala 66:21]
  assign _T_51 = rawA_sign == rawB_sign; // @[CompareRecFN.scala 72:34]
  assign _T_52 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62]
  assign _T_53 = _T_51 & _T_52; // @[CompareRecFN.scala 72:49]
  assign ordered_eq = bothZeros | _T_53; // @[CompareRecFN.scala 72:19]
  assign _T_56 = rawA_isNaN & ~rawA_sig[51]; // @[common.scala 81:46]
  assign _T_59 = rawB_isNaN & ~rawB_sig[51]; // @[common.scala 81:46]
  assign _T_60 = _T_56 | _T_59; // @[CompareRecFN.scala 75:32]
  assign invalid = _T_60 | ~ordered; // @[CompareRecFN.scala 75:58]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:11]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23]
endmodule
module ValExec_CompareRecF64_le(
  input         clock,
  input         reset,
  input  [63:0] io_a,
  input  [63:0] io_b,
  input         io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output        io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [64:0] compareRecFN_io_a; // @[ValExec_CompareRecFN.scala 94:30]
  wire [64:0] compareRecFN_io_b; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_lt; // @[ValExec_CompareRecFN.scala 94:30]
  wire  compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 94:30]
  wire [4:0] compareRecFN_io_exceptionFlags; // @[ValExec_CompareRecFN.scala 94:30]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_57; // @[Mux.scala 47:69]
  wire [5:0] _T_58; // @[Mux.scala 47:69]
  wire [5:0] _T_59; // @[Mux.scala 47:69]
  wire [5:0] _T_60; // @[Mux.scala 47:69]
  wire [5:0] _T_61; // @[Mux.scala 47:69]
  wire [5:0] _T_62; // @[Mux.scala 47:69]
  wire [5:0] _T_63; // @[Mux.scala 47:69]
  wire [5:0] _T_64; // @[Mux.scala 47:69]
  wire [5:0] _T_65; // @[Mux.scala 47:69]
  wire [5:0] _T_66; // @[Mux.scala 47:69]
  wire [5:0] _T_67; // @[Mux.scala 47:69]
  wire [5:0] _T_68; // @[Mux.scala 47:69]
  wire [5:0] _T_69; // @[Mux.scala 47:69]
  wire [5:0] _T_70; // @[Mux.scala 47:69]
  wire [5:0] _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [114:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_108; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_110; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_111; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_112; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_113; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_114; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_116; // @[rawFloatFromFN.scala 59:15]
  wire  _T_117; // @[rawFloatFromFN.scala 62:34]
  wire  _T_119; // @[rawFloatFromFN.scala 63:62]
  wire  _T_122; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_125; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_127; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_129; // @[Cat.scala 29:58]
  wire [2:0] _T_131; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_133; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_136; // @[Cat.scala 29:58]
  wire [3:0] _T_137; // @[Cat.scala 29:58]
  wire  _T_142; // @[rawFloatFromFN.scala 50:34]
  wire  _T_143; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_196; // @[Mux.scala 47:69]
  wire [5:0] _T_197; // @[Mux.scala 47:69]
  wire [5:0] _T_198; // @[Mux.scala 47:69]
  wire [5:0] _T_199; // @[Mux.scala 47:69]
  wire [5:0] _T_200; // @[Mux.scala 47:69]
  wire [5:0] _T_201; // @[Mux.scala 47:69]
  wire [5:0] _T_202; // @[Mux.scala 47:69]
  wire [5:0] _T_203; // @[Mux.scala 47:69]
  wire [5:0] _T_204; // @[Mux.scala 47:69]
  wire [5:0] _T_205; // @[Mux.scala 47:69]
  wire [5:0] _T_206; // @[Mux.scala 47:69]
  wire [5:0] _T_207; // @[Mux.scala 47:69]
  wire [5:0] _T_208; // @[Mux.scala 47:69]
  wire [5:0] _T_209; // @[Mux.scala 47:69]
  wire [5:0] _T_210; // @[Mux.scala 47:69]
  wire [5:0] _T_211; // @[Mux.scala 47:69]
  wire [5:0] _T_212; // @[Mux.scala 47:69]
  wire [5:0] _T_213; // @[Mux.scala 47:69]
  wire [5:0] _T_214; // @[Mux.scala 47:69]
  wire [5:0] _T_215; // @[Mux.scala 47:69]
  wire [5:0] _T_216; // @[Mux.scala 47:69]
  wire [5:0] _T_217; // @[Mux.scala 47:69]
  wire [5:0] _T_218; // @[Mux.scala 47:69]
  wire [5:0] _T_219; // @[Mux.scala 47:69]
  wire [5:0] _T_220; // @[Mux.scala 47:69]
  wire [5:0] _T_221; // @[Mux.scala 47:69]
  wire [5:0] _T_222; // @[Mux.scala 47:69]
  wire [5:0] _T_223; // @[Mux.scala 47:69]
  wire [5:0] _T_224; // @[Mux.scala 47:69]
  wire [5:0] _T_225; // @[Mux.scala 47:69]
  wire [5:0] _T_226; // @[Mux.scala 47:69]
  wire [5:0] _T_227; // @[Mux.scala 47:69]
  wire [5:0] _T_228; // @[Mux.scala 47:69]
  wire [5:0] _T_229; // @[Mux.scala 47:69]
  wire [5:0] _T_230; // @[Mux.scala 47:69]
  wire [5:0] _T_231; // @[Mux.scala 47:69]
  wire [5:0] _T_232; // @[Mux.scala 47:69]
  wire [5:0] _T_233; // @[Mux.scala 47:69]
  wire [5:0] _T_234; // @[Mux.scala 47:69]
  wire [5:0] _T_235; // @[Mux.scala 47:69]
  wire [5:0] _T_236; // @[Mux.scala 47:69]
  wire [5:0] _T_237; // @[Mux.scala 47:69]
  wire [5:0] _T_238; // @[Mux.scala 47:69]
  wire [5:0] _T_239; // @[Mux.scala 47:69]
  wire [5:0] _T_240; // @[Mux.scala 47:69]
  wire [5:0] _T_241; // @[Mux.scala 47:69]
  wire [5:0] _T_242; // @[Mux.scala 47:69]
  wire [5:0] _T_243; // @[Mux.scala 47:69]
  wire [5:0] _T_244; // @[Mux.scala 47:69]
  wire [5:0] _T_245; // @[Mux.scala 47:69]
  wire [5:0] _T_246; // @[Mux.scala 47:69]
  wire [114:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_247; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_249; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_250; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_251; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_252; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_253; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_255; // @[rawFloatFromFN.scala 59:15]
  wire  _T_256; // @[rawFloatFromFN.scala 62:34]
  wire  _T_258; // @[rawFloatFromFN.scala 63:62]
  wire  _T_261; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_264; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_266; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_268; // @[Cat.scala 29:58]
  wire [2:0] _T_270; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_272; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_275; // @[Cat.scala 29:58]
  wire [3:0] _T_276; // @[Cat.scala 29:58]
  wire  _T_279; // @[ValExec_CompareRecFN.scala 104:24]
  wire  _T_280; // @[ValExec_CompareRecFN.scala 105:35]
  CompareRecFN compareRecFN ( // @[ValExec_CompareRecFN.scala 94:30]
    .io_a(compareRecFN_io_a),
    .io_b(compareRecFN_io_b),
    .io_lt(compareRecFN_io_lt),
    .io_eq(compareRecFN_io_eq),
    .io_exceptionFlags(compareRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_a[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_a[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_57 = io_a[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_58 = io_a[2] ? 6'h31 : _T_57; // @[Mux.scala 47:69]
  assign _T_59 = io_a[3] ? 6'h30 : _T_58; // @[Mux.scala 47:69]
  assign _T_60 = io_a[4] ? 6'h2f : _T_59; // @[Mux.scala 47:69]
  assign _T_61 = io_a[5] ? 6'h2e : _T_60; // @[Mux.scala 47:69]
  assign _T_62 = io_a[6] ? 6'h2d : _T_61; // @[Mux.scala 47:69]
  assign _T_63 = io_a[7] ? 6'h2c : _T_62; // @[Mux.scala 47:69]
  assign _T_64 = io_a[8] ? 6'h2b : _T_63; // @[Mux.scala 47:69]
  assign _T_65 = io_a[9] ? 6'h2a : _T_64; // @[Mux.scala 47:69]
  assign _T_66 = io_a[10] ? 6'h29 : _T_65; // @[Mux.scala 47:69]
  assign _T_67 = io_a[11] ? 6'h28 : _T_66; // @[Mux.scala 47:69]
  assign _T_68 = io_a[12] ? 6'h27 : _T_67; // @[Mux.scala 47:69]
  assign _T_69 = io_a[13] ? 6'h26 : _T_68; // @[Mux.scala 47:69]
  assign _T_70 = io_a[14] ? 6'h25 : _T_69; // @[Mux.scala 47:69]
  assign _T_71 = io_a[15] ? 6'h24 : _T_70; // @[Mux.scala 47:69]
  assign _T_72 = io_a[16] ? 6'h23 : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = io_a[17] ? 6'h22 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = io_a[18] ? 6'h21 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = io_a[19] ? 6'h20 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = io_a[20] ? 6'h1f : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = io_a[21] ? 6'h1e : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = io_a[22] ? 6'h1d : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = io_a[23] ? 6'h1c : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = io_a[24] ? 6'h1b : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = io_a[25] ? 6'h1a : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = io_a[26] ? 6'h19 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = io_a[27] ? 6'h18 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = io_a[28] ? 6'h17 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = io_a[29] ? 6'h16 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = io_a[30] ? 6'h15 : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = io_a[31] ? 6'h14 : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = io_a[32] ? 6'h13 : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = io_a[33] ? 6'h12 : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = io_a[34] ? 6'h11 : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = io_a[35] ? 6'h10 : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = io_a[36] ? 6'hf : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = io_a[37] ? 6'he : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = io_a[38] ? 6'hd : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = io_a[39] ? 6'hc : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = io_a[40] ? 6'hb : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = io_a[41] ? 6'ha : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = io_a[42] ? 6'h9 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = io_a[43] ? 6'h8 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = io_a[44] ? 6'h7 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = io_a[45] ? 6'h6 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = io_a[46] ? 6'h5 : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = io_a[47] ? 6'h4 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = io_a[48] ? 6'h3 : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = io_a[49] ? 6'h2 : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = io_a[50] ? 6'h1 : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = io_a[51] ? 6'h0 : _T_106; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, io_a[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_108 = _GEN_0 << _T_107; // @[rawFloatFromFN.scala 54:36]
  assign _T_110 = {_T_108[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{6'd0}, _T_107}; // @[rawFloatFromFN.scala 57:26]
  assign _T_111 = _GEN_1 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_112 = _T_3 ? _T_111 : {{1'd0}, io_a[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_113 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{9'd0}, _T_113}; // @[rawFloatFromFN.scala 60:22]
  assign _T_114 = 11'h400 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_114}; // @[rawFloatFromFN.scala 59:15]
  assign _T_116 = _T_112 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_117 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_119 = _T_116[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_122 = _T_119 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_125 = {1'b0,$signed(_T_116)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_127 = _T_3 ? _T_110 : io_a[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_129 = {1'h0,~_T_117,_T_127}; // @[Cat.scala 29:58]
  assign _T_131 = _T_117 ? 3'h0 : _T_125[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_122}; // @[recFNFromFN.scala 48:79]
  assign _T_133 = _T_131 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_136 = {_T_125[8:0],_T_129[51:0]}; // @[Cat.scala 29:58]
  assign _T_137 = {io_a[63],_T_133}; // @[Cat.scala 29:58]
  assign _T_142 = io_b[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_143 = io_b[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_196 = io_b[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_197 = io_b[2] ? 6'h31 : _T_196; // @[Mux.scala 47:69]
  assign _T_198 = io_b[3] ? 6'h30 : _T_197; // @[Mux.scala 47:69]
  assign _T_199 = io_b[4] ? 6'h2f : _T_198; // @[Mux.scala 47:69]
  assign _T_200 = io_b[5] ? 6'h2e : _T_199; // @[Mux.scala 47:69]
  assign _T_201 = io_b[6] ? 6'h2d : _T_200; // @[Mux.scala 47:69]
  assign _T_202 = io_b[7] ? 6'h2c : _T_201; // @[Mux.scala 47:69]
  assign _T_203 = io_b[8] ? 6'h2b : _T_202; // @[Mux.scala 47:69]
  assign _T_204 = io_b[9] ? 6'h2a : _T_203; // @[Mux.scala 47:69]
  assign _T_205 = io_b[10] ? 6'h29 : _T_204; // @[Mux.scala 47:69]
  assign _T_206 = io_b[11] ? 6'h28 : _T_205; // @[Mux.scala 47:69]
  assign _T_207 = io_b[12] ? 6'h27 : _T_206; // @[Mux.scala 47:69]
  assign _T_208 = io_b[13] ? 6'h26 : _T_207; // @[Mux.scala 47:69]
  assign _T_209 = io_b[14] ? 6'h25 : _T_208; // @[Mux.scala 47:69]
  assign _T_210 = io_b[15] ? 6'h24 : _T_209; // @[Mux.scala 47:69]
  assign _T_211 = io_b[16] ? 6'h23 : _T_210; // @[Mux.scala 47:69]
  assign _T_212 = io_b[17] ? 6'h22 : _T_211; // @[Mux.scala 47:69]
  assign _T_213 = io_b[18] ? 6'h21 : _T_212; // @[Mux.scala 47:69]
  assign _T_214 = io_b[19] ? 6'h20 : _T_213; // @[Mux.scala 47:69]
  assign _T_215 = io_b[20] ? 6'h1f : _T_214; // @[Mux.scala 47:69]
  assign _T_216 = io_b[21] ? 6'h1e : _T_215; // @[Mux.scala 47:69]
  assign _T_217 = io_b[22] ? 6'h1d : _T_216; // @[Mux.scala 47:69]
  assign _T_218 = io_b[23] ? 6'h1c : _T_217; // @[Mux.scala 47:69]
  assign _T_219 = io_b[24] ? 6'h1b : _T_218; // @[Mux.scala 47:69]
  assign _T_220 = io_b[25] ? 6'h1a : _T_219; // @[Mux.scala 47:69]
  assign _T_221 = io_b[26] ? 6'h19 : _T_220; // @[Mux.scala 47:69]
  assign _T_222 = io_b[27] ? 6'h18 : _T_221; // @[Mux.scala 47:69]
  assign _T_223 = io_b[28] ? 6'h17 : _T_222; // @[Mux.scala 47:69]
  assign _T_224 = io_b[29] ? 6'h16 : _T_223; // @[Mux.scala 47:69]
  assign _T_225 = io_b[30] ? 6'h15 : _T_224; // @[Mux.scala 47:69]
  assign _T_226 = io_b[31] ? 6'h14 : _T_225; // @[Mux.scala 47:69]
  assign _T_227 = io_b[32] ? 6'h13 : _T_226; // @[Mux.scala 47:69]
  assign _T_228 = io_b[33] ? 6'h12 : _T_227; // @[Mux.scala 47:69]
  assign _T_229 = io_b[34] ? 6'h11 : _T_228; // @[Mux.scala 47:69]
  assign _T_230 = io_b[35] ? 6'h10 : _T_229; // @[Mux.scala 47:69]
  assign _T_231 = io_b[36] ? 6'hf : _T_230; // @[Mux.scala 47:69]
  assign _T_232 = io_b[37] ? 6'he : _T_231; // @[Mux.scala 47:69]
  assign _T_233 = io_b[38] ? 6'hd : _T_232; // @[Mux.scala 47:69]
  assign _T_234 = io_b[39] ? 6'hc : _T_233; // @[Mux.scala 47:69]
  assign _T_235 = io_b[40] ? 6'hb : _T_234; // @[Mux.scala 47:69]
  assign _T_236 = io_b[41] ? 6'ha : _T_235; // @[Mux.scala 47:69]
  assign _T_237 = io_b[42] ? 6'h9 : _T_236; // @[Mux.scala 47:69]
  assign _T_238 = io_b[43] ? 6'h8 : _T_237; // @[Mux.scala 47:69]
  assign _T_239 = io_b[44] ? 6'h7 : _T_238; // @[Mux.scala 47:69]
  assign _T_240 = io_b[45] ? 6'h6 : _T_239; // @[Mux.scala 47:69]
  assign _T_241 = io_b[46] ? 6'h5 : _T_240; // @[Mux.scala 47:69]
  assign _T_242 = io_b[47] ? 6'h4 : _T_241; // @[Mux.scala 47:69]
  assign _T_243 = io_b[48] ? 6'h3 : _T_242; // @[Mux.scala 47:69]
  assign _T_244 = io_b[49] ? 6'h2 : _T_243; // @[Mux.scala 47:69]
  assign _T_245 = io_b[50] ? 6'h1 : _T_244; // @[Mux.scala 47:69]
  assign _T_246 = io_b[51] ? 6'h0 : _T_245; // @[Mux.scala 47:69]
  assign _GEN_5 = {{63'd0}, io_b[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_247 = _GEN_5 << _T_246; // @[rawFloatFromFN.scala 54:36]
  assign _T_249 = {_T_247[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{6'd0}, _T_246}; // @[rawFloatFromFN.scala 57:26]
  assign _T_250 = _GEN_6 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_251 = _T_142 ? _T_250 : {{1'd0}, io_b[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_252 = _T_142 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{9'd0}, _T_252}; // @[rawFloatFromFN.scala 60:22]
  assign _T_253 = 11'h400 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_253}; // @[rawFloatFromFN.scala 59:15]
  assign _T_255 = _T_251 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_256 = _T_142 & _T_143; // @[rawFloatFromFN.scala 62:34]
  assign _T_258 = _T_255[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_261 = _T_258 & ~_T_143; // @[rawFloatFromFN.scala 66:33]
  assign _T_264 = {1'b0,$signed(_T_255)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_266 = _T_142 ? _T_249 : io_b[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_268 = {1'h0,~_T_256,_T_266}; // @[Cat.scala 29:58]
  assign _T_270 = _T_256 ? 3'h0 : _T_264[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_261}; // @[recFNFromFN.scala 48:79]
  assign _T_272 = _T_270 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_275 = {_T_264[8:0],_T_268[51:0]}; // @[Cat.scala 29:58]
  assign _T_276 = {io_b[63],_T_272}; // @[Cat.scala 29:58]
  assign _T_279 = io_actual_out == io_expected_out; // @[ValExec_CompareRecFN.scala 104:24]
  assign _T_280 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_CompareRecFN.scala 105:35]
  assign io_actual_out = compareRecFN_io_lt | compareRecFN_io_eq; // @[ValExec_CompareRecFN.scala 99:19]
  assign io_actual_exceptionFlags = compareRecFN_io_exceptionFlags; // @[ValExec_CompareRecFN.scala 100:30]
  assign io_check = 1'h1; // @[ValExec_CompareRecFN.scala 102:14]
  assign io_pass = _T_279 & _T_280; // @[ValExec_CompareRecFN.scala 103:13]
  assign compareRecFN_io_a = {_T_137,_T_136}; // @[ValExec_CompareRecFN.scala 95:23]
  assign compareRecFN_io_b = {_T_276,_T_275}; // @[ValExec_CompareRecFN.scala 96:23]
endmodule
