module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [53:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [16:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [13:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 108:24]
  wire  _T_5; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [13:0] adjustedSig; // @[Cat.scala 29:58]
  wire [64:0] _T_8; // @[primitives.scala 77:58]
  wire [7:0] _T_14; // @[Bitwise.scala 102:31]
  wire [7:0] _T_16; // @[Bitwise.scala 102:65]
  wire [7:0] _T_18; // @[Bitwise.scala 102:75]
  wire [7:0] _T_19; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_0; // @[Bitwise.scala 102:31]
  wire [7:0] _T_24; // @[Bitwise.scala 102:31]
  wire [7:0] _T_26; // @[Bitwise.scala 102:65]
  wire [7:0] _T_28; // @[Bitwise.scala 102:75]
  wire [7:0] _T_29; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [7:0] _T_34; // @[Bitwise.scala 102:31]
  wire [7:0] _T_36; // @[Bitwise.scala 102:65]
  wire [7:0] _T_38; // @[Bitwise.scala 102:75]
  wire [7:0] _T_39; // @[Bitwise.scala 102:39]
  wire [13:0] _T_52; // @[Cat.scala 29:58]
  wire [13:0] _T_54; // @[Cat.scala 29:58]
  wire [13:0] _T_56; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [13:0] _T_57; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_58; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [13:0] _T_59; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_60; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_61; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_62; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_63; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_64; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_65; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [13:0] _T_66; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [12:0] _T_68; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_69; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_71; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [12:0] _T_73; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [12:0] _T_75; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [13:0] _T_77; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_79; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [12:0] _T_81; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [12:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] _T_82; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] _T_83; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_85; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [13:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [14:0] _T_86; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [5:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [9:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [10:0] _T_91; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_100; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_103; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_104; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_105; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire [8:0] _T_109; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_110; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_111; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_115; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_121; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_122; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_123; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_124; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_126; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _T_131; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_133; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_135; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_136; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_138; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_139; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [5:0] _T_140; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [5:0] _T_142; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [5:0] _T_144; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [5:0] _T_146; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [5:0] _T_147; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [5:0] _T_149; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [5:0] _T_150; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [5:0] _T_152; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [5:0] _T_153; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [5:0] _T_154; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [5:0] _T_155; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [5:0] _T_156; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [5:0] _T_157; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [5:0] _T_158; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [5:0] _T_159; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [5:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_160; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [9:0] _T_162; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [9:0] _T_163; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] _T_165; // @[Bitwise.scala 71:12]
  wire [9:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [6:0] _T_166; // @[Cat.scala 29:58]
  wire [1:0] _T_168; // @[Cat.scala 29:58]
  wire [2:0] _T_170; // @[Cat.scala 29:58]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign sAdjustedExp = $signed(io_in_sExp) - 13'sh7e0; // @[RoundAnyRawFNToRecFN.scala 108:24]
  assign _T_5 = io_in_sig[40:0] != 41'h0; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[53:41],_T_5}; // @[Cat.scala 29:58]
  assign _T_8 = -65'sh10000000000000000 >>> ~sAdjustedExp[5:0]; // @[primitives.scala 77:58]
  assign _T_14 = {{4'd0}, _T_8[14:11]}; // @[Bitwise.scala 102:31]
  assign _T_16 = {_T_8[10:7], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_18 = _T_16 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_19 = _T_14 | _T_18; // @[Bitwise.scala 102:39]
  assign _GEN_0 = {{2'd0}, _T_19[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_24 = _GEN_0 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_26 = {_T_19[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_28 = _T_26 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_29 = _T_24 | _T_28; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{1'd0}, _T_29[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_34 = _GEN_1 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_36 = {_T_29[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_38 = _T_36 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_39 = _T_34 | _T_38; // @[Bitwise.scala 102:39]
  assign _T_52 = {_T_39,_T_8[15],_T_8[16],_T_8[17],_T_8[18],2'h3}; // @[Cat.scala 29:58]
  assign _T_54 = {1'h0,_T_52[13:1]}; // @[Cat.scala 29:58]
  assign _T_56 = ~_T_54 & _T_52; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_57 = adjustedSig & _T_56; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_58 = _T_57 != 14'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_59 = adjustedSig & _T_54; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_60 = _T_59 != 14'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_61 = _T_58 | _T_60; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_62 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_63 = _T_62 & _T_58; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_64 = roundMagUp & _T_61; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_65 = _T_63 | _T_64; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_66 = adjustedSig | _T_52; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_68 = _T_66[13:2] + 12'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_69 = roundingMode_near_even & _T_58; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_71 = _T_69 & ~_T_60; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_73 = _T_71 ? _T_52[13:1] : 13'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_75 = _T_68 & ~_T_73; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_77 = adjustedSig & ~_T_52; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_79 = roundingMode_odd & _T_61; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_81 = _T_79 ? _T_56[13:1] : 13'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_2 = {{1'd0}, _T_77[13:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_82 = _GEN_2 | _T_81; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_83 = _T_65 ? _T_75 : _T_82; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_85 = {1'b0,$signed(_T_83[12:11])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_3 = {{11{_T_85[2]}},_T_85}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_86 = $signed(sAdjustedExp) + $signed(_GEN_3); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_86[5:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_83[9:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign _T_91 = _T_86[14:4]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_91) >= 11'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_86) < 15'sh8; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_100 = adjustedSig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_103 = _T_62 & adjustedSig[1]; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_104 = roundMagUp & _T_100; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_105 = _T_103 | _T_104; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_109 = sAdjustedExp[13:5]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_110 = $signed(_T_109) <= 9'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_111 = _T_61 & _T_110; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_115 = _T_111 & _T_52[2]; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_121 = io_detectTininess & ~_T_52[3]; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_122 = _T_121 & _T_83[11]; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_123 = _T_122 & _T_58; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_124 = _T_123 & _T_105; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_126 = _T_115 & ~_T_124; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_126; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_61; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign _T_131 = ~isNaNOut & ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_131 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_133 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_133; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_62 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_135 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_136 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_135 & _T_136; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_138 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = io_in_isInf | _T_138; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_139 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_140 = _T_139 ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_142 = common_expOut & ~_T_140; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_144 = pegMinNonzeroMagOut ? 6'h37 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_146 = _T_142 & ~_T_144; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_147 = pegMaxFiniteMagOut ? 6'h10 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_149 = _T_146 & ~_T_147; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_150 = notNaN_isInfOut ? 6'h8 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_152 = _T_149 & ~_T_150; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_153 = pegMinNonzeroMagOut ? 6'h8 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_154 = _T_152 | _T_153; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_155 = pegMaxFiniteMagOut ? 6'h2f : 6'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_156 = _T_154 | _T_155; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_157 = notNaN_isInfOut ? 6'h30 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_158 = _T_156 | _T_157; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_159 = isNaNOut ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_158 | _T_159; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_160 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_161 = _T_160 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_162 = isNaNOut ? 10'h200 : 10'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_163 = _T_161 ? _T_162 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_165 = pegMaxFiniteMagOut ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign fractOut = _T_163 | _T_165; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_166 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_168 = {underflow,inexact}; // @[Cat.scala 29:58]
  assign _T_170 = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_166,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_170,_T_168}; // @[RoundAnyRawFNToRecFN.scala 285:23]
endmodule
module RecFNToRecFN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [16:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  RoundAnyRawFNToRecFN_io_invalidExc; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isNaN; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isInf; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_isZero; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_in_sign; // @[RecFNToRecFN.scala 72:19]
  wire [12:0] RoundAnyRawFNToRecFN_io_in_sExp; // @[RecFNToRecFN.scala 72:19]
  wire [53:0] RoundAnyRawFNToRecFN_io_in_sig; // @[RecFNToRecFN.scala 72:19]
  wire [2:0] RoundAnyRawFNToRecFN_io_roundingMode; // @[RecFNToRecFN.scala 72:19]
  wire  RoundAnyRawFNToRecFN_io_detectTininess; // @[RecFNToRecFN.scala 72:19]
  wire [16:0] RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 72:19]
  wire [4:0] RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 72:19]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [53:0] rawIn_sig; // @[Cat.scala 29:58]
  RoundAnyRawFNToRecFN RoundAnyRawFNToRecFN ( // @[RecFNToRecFN.scala 72:19]
    .io_invalidExc(RoundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(RoundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(RoundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(RoundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(RoundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(RoundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(RoundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(RoundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(RoundAnyRawFNToRecFN_io_detectTininess),
    .io_out(RoundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(RoundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn_isNaN = _T_4 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  assign _T_14 = {1'h0,~rawIn_isZero}; // @[Cat.scala 29:58]
  assign rawIn_sig = {1'h0,~rawIn_isZero,io_in[51:0]}; // @[Cat.scala 29:58]
  assign io_out = RoundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 85:27]
  assign io_exceptionFlags = RoundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 86:27]
  assign RoundAnyRawFNToRecFN_io_invalidExc = rawIn_isNaN & ~rawIn_sig[51]; // @[RecFNToRecFN.scala 80:48]
  assign RoundAnyRawFNToRecFN_io_in_isNaN = _T_4 & io_in[61]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isInf = _T_4 & ~io_in[61]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_isZero = io_in[63:61] == 3'h0; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sign = io_in[64]; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(io_in[63:52])}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_in_sig = {_T_14,io_in[51:0]}; // @[RecFNToRecFN.scala 82:48]
  assign RoundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RecFNToRecFN.scala 83:48]
  assign RoundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RecFNToRecFN.scala 84:48]
endmodule
module ValExec_RecF64ToRecF16(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [15:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [16:0] io_expected_recOut,
  output [16:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [64:0] recFNToRecFN_io_in; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire [2:0] recFNToRecFN_io_roundingMode; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire  recFNToRecFN_io_detectTininess; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire [16:0] recFNToRecFN_io_out; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire [4:0] recFNToRecFN_io_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 68:15]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_57; // @[Mux.scala 47:69]
  wire [5:0] _T_58; // @[Mux.scala 47:69]
  wire [5:0] _T_59; // @[Mux.scala 47:69]
  wire [5:0] _T_60; // @[Mux.scala 47:69]
  wire [5:0] _T_61; // @[Mux.scala 47:69]
  wire [5:0] _T_62; // @[Mux.scala 47:69]
  wire [5:0] _T_63; // @[Mux.scala 47:69]
  wire [5:0] _T_64; // @[Mux.scala 47:69]
  wire [5:0] _T_65; // @[Mux.scala 47:69]
  wire [5:0] _T_66; // @[Mux.scala 47:69]
  wire [5:0] _T_67; // @[Mux.scala 47:69]
  wire [5:0] _T_68; // @[Mux.scala 47:69]
  wire [5:0] _T_69; // @[Mux.scala 47:69]
  wire [5:0] _T_70; // @[Mux.scala 47:69]
  wire [5:0] _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [114:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_108; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_110; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_111; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_112; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_113; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_114; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_116; // @[rawFloatFromFN.scala 59:15]
  wire  _T_117; // @[rawFloatFromFN.scala 62:34]
  wire  _T_119; // @[rawFloatFromFN.scala 63:62]
  wire  _T_122; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_125; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_127; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_129; // @[Cat.scala 29:58]
  wire [2:0] _T_131; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_133; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_136; // @[Cat.scala 29:58]
  wire [3:0] _T_137; // @[Cat.scala 29:58]
  wire  _T_142; // @[rawFloatFromFN.scala 50:34]
  wire  _T_143; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_154; // @[Mux.scala 47:69]
  wire [3:0] _T_155; // @[Mux.scala 47:69]
  wire [3:0] _T_156; // @[Mux.scala 47:69]
  wire [3:0] _T_157; // @[Mux.scala 47:69]
  wire [3:0] _T_158; // @[Mux.scala 47:69]
  wire [3:0] _T_159; // @[Mux.scala 47:69]
  wire [3:0] _T_160; // @[Mux.scala 47:69]
  wire [3:0] _T_161; // @[Mux.scala 47:69]
  wire [3:0] _T_162; // @[Mux.scala 47:69]
  wire [24:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_163; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_165; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_166; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_167; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_168; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_169; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_171; // @[rawFloatFromFN.scala 59:15]
  wire  _T_172; // @[rawFloatFromFN.scala 62:34]
  wire  _T_174; // @[rawFloatFromFN.scala 63:62]
  wire  _T_177; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_180; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_182; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_184; // @[Cat.scala 29:58]
  wire [2:0] _T_186; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_188; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_191; // @[Cat.scala 29:58]
  wire [3:0] _T_192; // @[Cat.scala 29:58]
  wire  _T_197; // @[tests.scala 48:26]
  wire  _T_199; // @[tests.scala 48:55]
  wire  _T_200; // @[tests.scala 48:39]
  wire  _T_201; // @[tests.scala 49:20]
  wire  _T_204; // @[tests.scala 49:54]
  wire  _T_205; // @[tests.scala 49:31]
  wire  _T_207; // @[tests.scala 50:30]
  wire  _T_209; // @[tests.scala 50:66]
  wire  _T_210; // @[tests.scala 50:16]
  wire  _T_211; // @[tests.scala 48:12]
  wire  _T_212; // @[ValExec_RecFNToRecFN.scala 84:35]
  RecFNToRecFN recFNToRecFN ( // @[ValExec_RecFNToRecFN.scala 68:15]
    .io_in(recFNToRecFN_io_in),
    .io_roundingMode(recFNToRecFN_io_roundingMode),
    .io_detectTininess(recFNToRecFN_io_detectTininess),
    .io_out(recFNToRecFN_io_out),
    .io_exceptionFlags(recFNToRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_in[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_in[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_57 = io_in[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_58 = io_in[2] ? 6'h31 : _T_57; // @[Mux.scala 47:69]
  assign _T_59 = io_in[3] ? 6'h30 : _T_58; // @[Mux.scala 47:69]
  assign _T_60 = io_in[4] ? 6'h2f : _T_59; // @[Mux.scala 47:69]
  assign _T_61 = io_in[5] ? 6'h2e : _T_60; // @[Mux.scala 47:69]
  assign _T_62 = io_in[6] ? 6'h2d : _T_61; // @[Mux.scala 47:69]
  assign _T_63 = io_in[7] ? 6'h2c : _T_62; // @[Mux.scala 47:69]
  assign _T_64 = io_in[8] ? 6'h2b : _T_63; // @[Mux.scala 47:69]
  assign _T_65 = io_in[9] ? 6'h2a : _T_64; // @[Mux.scala 47:69]
  assign _T_66 = io_in[10] ? 6'h29 : _T_65; // @[Mux.scala 47:69]
  assign _T_67 = io_in[11] ? 6'h28 : _T_66; // @[Mux.scala 47:69]
  assign _T_68 = io_in[12] ? 6'h27 : _T_67; // @[Mux.scala 47:69]
  assign _T_69 = io_in[13] ? 6'h26 : _T_68; // @[Mux.scala 47:69]
  assign _T_70 = io_in[14] ? 6'h25 : _T_69; // @[Mux.scala 47:69]
  assign _T_71 = io_in[15] ? 6'h24 : _T_70; // @[Mux.scala 47:69]
  assign _T_72 = io_in[16] ? 6'h23 : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = io_in[17] ? 6'h22 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = io_in[18] ? 6'h21 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = io_in[19] ? 6'h20 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = io_in[20] ? 6'h1f : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = io_in[21] ? 6'h1e : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = io_in[22] ? 6'h1d : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = io_in[23] ? 6'h1c : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = io_in[24] ? 6'h1b : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = io_in[25] ? 6'h1a : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = io_in[26] ? 6'h19 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = io_in[27] ? 6'h18 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = io_in[28] ? 6'h17 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = io_in[29] ? 6'h16 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = io_in[30] ? 6'h15 : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = io_in[31] ? 6'h14 : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = io_in[32] ? 6'h13 : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = io_in[33] ? 6'h12 : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = io_in[34] ? 6'h11 : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = io_in[35] ? 6'h10 : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = io_in[36] ? 6'hf : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = io_in[37] ? 6'he : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = io_in[38] ? 6'hd : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = io_in[39] ? 6'hc : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = io_in[40] ? 6'hb : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = io_in[41] ? 6'ha : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = io_in[42] ? 6'h9 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = io_in[43] ? 6'h8 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = io_in[44] ? 6'h7 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = io_in[45] ? 6'h6 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = io_in[46] ? 6'h5 : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = io_in[47] ? 6'h4 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = io_in[48] ? 6'h3 : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = io_in[49] ? 6'h2 : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = io_in[50] ? 6'h1 : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = io_in[51] ? 6'h0 : _T_106; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, io_in[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_108 = _GEN_0 << _T_107; // @[rawFloatFromFN.scala 54:36]
  assign _T_110 = {_T_108[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{6'd0}, _T_107}; // @[rawFloatFromFN.scala 57:26]
  assign _T_111 = _GEN_1 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_112 = _T_3 ? _T_111 : {{1'd0}, io_in[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_113 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{9'd0}, _T_113}; // @[rawFloatFromFN.scala 60:22]
  assign _T_114 = 11'h400 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_114}; // @[rawFloatFromFN.scala 59:15]
  assign _T_116 = _T_112 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_117 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_119 = _T_116[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_122 = _T_119 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_125 = {1'b0,$signed(_T_116)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_127 = _T_3 ? _T_110 : io_in[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_129 = {1'h0,~_T_117,_T_127}; // @[Cat.scala 29:58]
  assign _T_131 = _T_117 ? 3'h0 : _T_125[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_122}; // @[recFNFromFN.scala 48:79]
  assign _T_133 = _T_131 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_136 = {_T_125[8:0],_T_129[51:0]}; // @[Cat.scala 29:58]
  assign _T_137 = {io_in[63],_T_133}; // @[Cat.scala 29:58]
  assign _T_142 = io_expected_out[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_143 = io_expected_out[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_154 = io_expected_out[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_155 = io_expected_out[2] ? 4'h7 : _T_154; // @[Mux.scala 47:69]
  assign _T_156 = io_expected_out[3] ? 4'h6 : _T_155; // @[Mux.scala 47:69]
  assign _T_157 = io_expected_out[4] ? 4'h5 : _T_156; // @[Mux.scala 47:69]
  assign _T_158 = io_expected_out[5] ? 4'h4 : _T_157; // @[Mux.scala 47:69]
  assign _T_159 = io_expected_out[6] ? 4'h3 : _T_158; // @[Mux.scala 47:69]
  assign _T_160 = io_expected_out[7] ? 4'h2 : _T_159; // @[Mux.scala 47:69]
  assign _T_161 = io_expected_out[8] ? 4'h1 : _T_160; // @[Mux.scala 47:69]
  assign _T_162 = io_expected_out[9] ? 4'h0 : _T_161; // @[Mux.scala 47:69]
  assign _GEN_5 = {{15'd0}, io_expected_out[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_163 = _GEN_5 << _T_162; // @[rawFloatFromFN.scala 54:36]
  assign _T_165 = {_T_163[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{2'd0}, _T_162}; // @[rawFloatFromFN.scala 57:26]
  assign _T_166 = _GEN_6 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_167 = _T_142 ? _T_166 : {{1'd0}, io_expected_out[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_168 = _T_142 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{3'd0}, _T_168}; // @[rawFloatFromFN.scala 60:22]
  assign _T_169 = 5'h10 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_169}; // @[rawFloatFromFN.scala 59:15]
  assign _T_171 = _T_167 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_172 = _T_142 & _T_143; // @[rawFloatFromFN.scala 62:34]
  assign _T_174 = _T_171[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_177 = _T_174 & ~_T_143; // @[rawFloatFromFN.scala 66:33]
  assign _T_180 = {1'b0,$signed(_T_171)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_182 = _T_142 ? _T_165 : io_expected_out[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_184 = {1'h0,~_T_172,_T_182}; // @[Cat.scala 29:58]
  assign _T_186 = _T_172 ? 3'h0 : _T_180[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_177}; // @[recFNFromFN.scala 48:79]
  assign _T_188 = _T_186 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_191 = {_T_180[2:0],_T_184[9:0]}; // @[Cat.scala 29:58]
  assign _T_192 = {io_expected_out[15],_T_188}; // @[Cat.scala 29:58]
  assign _T_197 = io_actual_out[15:13] == 3'h0; // @[tests.scala 48:26]
  assign _T_199 = io_actual_out[15:13] == 3'h7; // @[tests.scala 48:55]
  assign _T_200 = _T_197 | _T_199; // @[tests.scala 48:39]
  assign _T_201 = io_actual_out[16:13] == io_expected_recOut[16:13]; // @[tests.scala 49:20]
  assign _T_204 = io_actual_out[9:0] == io_expected_recOut[9:0]; // @[tests.scala 49:54]
  assign _T_205 = _T_201 & _T_204; // @[tests.scala 49:31]
  assign _T_207 = io_actual_out[15:13] == 3'h6; // @[tests.scala 50:30]
  assign _T_209 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_210 = _T_207 ? _T_201 : _T_209; // @[tests.scala 50:16]
  assign _T_211 = _T_200 ? _T_205 : _T_210; // @[tests.scala 48:12]
  assign _T_212 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 84:35]
  assign io_expected_recOut = {_T_192,_T_191}; // @[ValExec_RecFNToRecFN.scala 74:24]
  assign io_actual_out = recFNToRecFN_io_out; // @[ValExec_RecFNToRecFN.scala 77:19]
  assign io_actual_exceptionFlags = recFNToRecFN_io_exceptionFlags; // @[ValExec_RecFNToRecFN.scala 78:30]
  assign io_check = 1'h1; // @[ValExec_RecFNToRecFN.scala 80:14]
  assign io_pass = _T_211 & _T_212; // @[ValExec_RecFNToRecFN.scala 81:13]
  assign recFNToRecFN_io_in = {_T_137,_T_136}; // @[ValExec_RecFNToRecFN.scala 70:24]
  assign recFNToRecFN_io_roundingMode = io_roundingMode; // @[ValExec_RecFNToRecFN.scala 71:36]
  assign recFNToRecFN_io_detectTininess = io_detectTininess; // @[ValExec_RecFNToRecFN.scala 72:36]
endmodule
