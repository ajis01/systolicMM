module MixedVecConnectWithSeqTester(
  input   clock,
  input   reset
);
  wire  _T_13; // @[MixedVecSpec.scala 138:7]
  assign _T_13 = reset == 1'h0; // @[MixedVecSpec.scala 138:7]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $finish; // @[MixedVecSpec.scala 138:7]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
