module RoundAnyRawFNToRecFN(
  input         io_in_isZero,
  input  [7:0]  io_in_sExp,
  input  [32:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [16:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire [8:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 108:24]
  wire  _T_5; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [13:0] adjustedSig; // @[Cat.scala 29:58]
  wire [13:0] _T_12; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_13; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [13:0] _T_14; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_15; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_17; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_18; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_19; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_20; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [13:0] _T_21; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [12:0] _T_23; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_24; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_26; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [12:0] _T_28; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [12:0] _T_30; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [13:0] _T_32; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_34; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [12:0] _T_36; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [12:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] _T_37; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] _T_38; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [8:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [9:0] _T_41; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [5:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [9:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [5:0] _T_46; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  _T_68; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire [5:0] _T_75; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [5:0] _T_77; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [5:0] _T_82; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [5:0] _T_84; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [5:0] _T_85; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [5:0] _T_87; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [5:0] _T_90; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [5:0] _T_91; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [5:0] _T_92; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [5:0] expOut; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [9:0] _T_98; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] _T_100; // @[Bitwise.scala 71:12]
  wire [9:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [6:0] _T_101; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[Cat.scala 29:58]
  wire [2:0] _T_105; // @[Cat.scala 29:58]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign sAdjustedExp = $signed(io_in_sExp) - 8'sh20; // @[RoundAnyRawFNToRecFN.scala 108:24]
  assign _T_5 = io_in_sig[19:0] != 20'h0; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {io_in_sig[32:20],_T_5}; // @[Cat.scala 29:58]
  assign _T_12 = adjustedSig & 14'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_13 = _T_12 != 14'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_14 = adjustedSig & 14'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_15 = _T_14 != 14'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign common_inexact = _T_13 | _T_15; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_17 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_18 = _T_17 & _T_13; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_19 = roundingMode_max & common_inexact; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_20 = _T_18 | _T_19; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_21 = adjustedSig | 14'h3; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_23 = _T_21[13:2] + 12'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_24 = roundingMode_near_even & _T_13; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_26 = _T_24 & ~_T_15; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_28 = _T_26 ? 13'h1 : 13'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_30 = _T_23 & ~_T_28; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_32 = adjustedSig & 14'h3ffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_34 = roundingMode_odd & common_inexact; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_36 = _T_34 ? 13'h1 : 13'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_0 = {{1'd0}, _T_32[13:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_37 = _GEN_0 | _T_36; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_38 = _T_20 ? _T_30 : _T_37; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_40 = {1'b0,$signed(_T_38[12:11])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_1 = {{6{_T_40[2]}},_T_40}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_41 = $signed(sAdjustedExp) + $signed(_GEN_1); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_41[5:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = _T_38[9:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign _T_46 = _T_41[9:4]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_46) >= 6'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign _T_68 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_68; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_17 | roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign notNaN_isInfOut = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign _T_75 = io_in_isZero ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_77 = common_expOut & ~_T_75; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_82 = pegMaxFiniteMagOut ? 6'h10 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_84 = _T_77 & ~_T_82; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_85 = notNaN_isInfOut ? 6'h8 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_87 = _T_84 & ~_T_85; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_90 = pegMaxFiniteMagOut ? 6'h2f : 6'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_91 = _T_87 | _T_90; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_92 = notNaN_isInfOut ? 6'h30 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign expOut = _T_91 | _T_92; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_98 = io_in_isZero ? 10'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_100 = pegMaxFiniteMagOut ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign fractOut = _T_98 | _T_100; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_101 = {1'h0,expOut}; // @[Cat.scala 29:58]
  assign _T_103 = {1'h0,inexact}; // @[Cat.scala 29:58]
  assign _T_105 = {2'h0,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_101,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_105,_T_103}; // @[RoundAnyRawFNToRecFN.scala 285:23]
endmodule
module INToRecFN(
  input  [31:0] io_in,
  input  [2:0]  io_roundingMode,
  output [16:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire [7:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [32:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15]
  wire [16:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15]
  wire [63:0] _T_5; // @[Cat.scala 29:58]
  wire [4:0] _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_48; // @[Mux.scala 47:69]
  wire [4:0] _T_49; // @[Mux.scala 47:69]
  wire [4:0] _T_50; // @[Mux.scala 47:69]
  wire [4:0] _T_51; // @[Mux.scala 47:69]
  wire [4:0] _T_52; // @[Mux.scala 47:69]
  wire [4:0] _T_53; // @[Mux.scala 47:69]
  wire [4:0] _T_54; // @[Mux.scala 47:69]
  wire [4:0] _T_55; // @[Mux.scala 47:69]
  wire [4:0] _T_56; // @[Mux.scala 47:69]
  wire [4:0] _T_57; // @[Mux.scala 47:69]
  wire [4:0] _T_58; // @[Mux.scala 47:69]
  wire [4:0] _T_59; // @[Mux.scala 47:69]
  wire [4:0] _T_60; // @[Mux.scala 47:69]
  wire [4:0] _T_61; // @[Mux.scala 47:69]
  wire [4:0] _T_62; // @[Mux.scala 47:69]
  wire [4:0] _T_63; // @[Mux.scala 47:69]
  wire [4:0] _T_64; // @[Mux.scala 47:69]
  wire [4:0] _T_65; // @[Mux.scala 47:69]
  wire [4:0] _T_66; // @[Mux.scala 47:69]
  wire [4:0] _T_67; // @[Mux.scala 47:69]
  wire [4:0] _T_68; // @[Mux.scala 47:69]
  wire [4:0] _T_69; // @[Mux.scala 47:69]
  wire [62:0] _GEN_0; // @[rawFloatFromIN.scala 55:22]
  wire [62:0] _T_70; // @[rawFloatFromIN.scala 55:22]
  wire [6:0] _T_76; // @[Cat.scala 29:58]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign _T_5 = {32'h0,io_in}; // @[Cat.scala 29:58]
  assign _T_39 = _T_5[1] ? 5'h1e : 5'h1f; // @[Mux.scala 47:69]
  assign _T_40 = _T_5[2] ? 5'h1d : _T_39; // @[Mux.scala 47:69]
  assign _T_41 = _T_5[3] ? 5'h1c : _T_40; // @[Mux.scala 47:69]
  assign _T_42 = _T_5[4] ? 5'h1b : _T_41; // @[Mux.scala 47:69]
  assign _T_43 = _T_5[5] ? 5'h1a : _T_42; // @[Mux.scala 47:69]
  assign _T_44 = _T_5[6] ? 5'h19 : _T_43; // @[Mux.scala 47:69]
  assign _T_45 = _T_5[7] ? 5'h18 : _T_44; // @[Mux.scala 47:69]
  assign _T_46 = _T_5[8] ? 5'h17 : _T_45; // @[Mux.scala 47:69]
  assign _T_47 = _T_5[9] ? 5'h16 : _T_46; // @[Mux.scala 47:69]
  assign _T_48 = _T_5[10] ? 5'h15 : _T_47; // @[Mux.scala 47:69]
  assign _T_49 = _T_5[11] ? 5'h14 : _T_48; // @[Mux.scala 47:69]
  assign _T_50 = _T_5[12] ? 5'h13 : _T_49; // @[Mux.scala 47:69]
  assign _T_51 = _T_5[13] ? 5'h12 : _T_50; // @[Mux.scala 47:69]
  assign _T_52 = _T_5[14] ? 5'h11 : _T_51; // @[Mux.scala 47:69]
  assign _T_53 = _T_5[15] ? 5'h10 : _T_52; // @[Mux.scala 47:69]
  assign _T_54 = _T_5[16] ? 5'hf : _T_53; // @[Mux.scala 47:69]
  assign _T_55 = _T_5[17] ? 5'he : _T_54; // @[Mux.scala 47:69]
  assign _T_56 = _T_5[18] ? 5'hd : _T_55; // @[Mux.scala 47:69]
  assign _T_57 = _T_5[19] ? 5'hc : _T_56; // @[Mux.scala 47:69]
  assign _T_58 = _T_5[20] ? 5'hb : _T_57; // @[Mux.scala 47:69]
  assign _T_59 = _T_5[21] ? 5'ha : _T_58; // @[Mux.scala 47:69]
  assign _T_60 = _T_5[22] ? 5'h9 : _T_59; // @[Mux.scala 47:69]
  assign _T_61 = _T_5[23] ? 5'h8 : _T_60; // @[Mux.scala 47:69]
  assign _T_62 = _T_5[24] ? 5'h7 : _T_61; // @[Mux.scala 47:69]
  assign _T_63 = _T_5[25] ? 5'h6 : _T_62; // @[Mux.scala 47:69]
  assign _T_64 = _T_5[26] ? 5'h5 : _T_63; // @[Mux.scala 47:69]
  assign _T_65 = _T_5[27] ? 5'h4 : _T_64; // @[Mux.scala 47:69]
  assign _T_66 = _T_5[28] ? 5'h3 : _T_65; // @[Mux.scala 47:69]
  assign _T_67 = _T_5[29] ? 5'h2 : _T_66; // @[Mux.scala 47:69]
  assign _T_68 = _T_5[30] ? 5'h1 : _T_67; // @[Mux.scala 47:69]
  assign _T_69 = _T_5[31] ? 5'h0 : _T_68; // @[Mux.scala 47:69]
  assign _GEN_0 = {{31'd0}, _T_5[31:0]}; // @[rawFloatFromIN.scala 55:22]
  assign _T_70 = _GEN_0 << _T_69; // @[rawFloatFromIN.scala 55:22]
  assign _T_76 = {2'h2,~_T_69}; // @[Cat.scala 29:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_70[31]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_76)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_70[31:0]}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44]
endmodule
module ValExec_UI32ToRecF16(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [15:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [16:0] io_expected_recOut,
  output [16:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [31:0] iNToRecFN_io_in; // @[ValExec_INToRecFN.scala 66:27]
  wire [2:0] iNToRecFN_io_roundingMode; // @[ValExec_INToRecFN.scala 66:27]
  wire [16:0] iNToRecFN_io_out; // @[ValExec_INToRecFN.scala 66:27]
  wire [4:0] iNToRecFN_io_exceptionFlags; // @[ValExec_INToRecFN.scala 66:27]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_15; // @[Mux.scala 47:69]
  wire [3:0] _T_16; // @[Mux.scala 47:69]
  wire [3:0] _T_17; // @[Mux.scala 47:69]
  wire [3:0] _T_18; // @[Mux.scala 47:69]
  wire [3:0] _T_19; // @[Mux.scala 47:69]
  wire [3:0] _T_20; // @[Mux.scala 47:69]
  wire [3:0] _T_21; // @[Mux.scala 47:69]
  wire [3:0] _T_22; // @[Mux.scala 47:69]
  wire [3:0] _T_23; // @[Mux.scala 47:69]
  wire [24:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_24; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_26; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_27; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_28; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_29; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_30; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_32; // @[rawFloatFromFN.scala 59:15]
  wire  _T_33; // @[rawFloatFromFN.scala 62:34]
  wire  _T_35; // @[rawFloatFromFN.scala 63:62]
  wire  _T_38; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_41; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_43; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_45; // @[Cat.scala 29:58]
  wire [2:0] _T_47; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_49; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_52; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[Cat.scala 29:58]
  wire  _T_58; // @[tests.scala 48:26]
  wire  _T_60; // @[tests.scala 48:55]
  wire  _T_61; // @[tests.scala 48:39]
  wire  _T_62; // @[tests.scala 49:20]
  wire  _T_65; // @[tests.scala 49:54]
  wire  _T_66; // @[tests.scala 49:31]
  wire  _T_68; // @[tests.scala 50:30]
  wire  _T_70; // @[tests.scala 50:66]
  wire  _T_71; // @[tests.scala 50:16]
  wire  _T_72; // @[tests.scala 48:12]
  wire  _T_73; // @[ValExec_INToRecFN.scala 80:35]
  INToRecFN iNToRecFN ( // @[ValExec_INToRecFN.scala 66:27]
    .io_in(iNToRecFN_io_in),
    .io_roundingMode(iNToRecFN_io_roundingMode),
    .io_out(iNToRecFN_io_out),
    .io_exceptionFlags(iNToRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_expected_out[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_expected_out[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_15 = io_expected_out[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_16 = io_expected_out[2] ? 4'h7 : _T_15; // @[Mux.scala 47:69]
  assign _T_17 = io_expected_out[3] ? 4'h6 : _T_16; // @[Mux.scala 47:69]
  assign _T_18 = io_expected_out[4] ? 4'h5 : _T_17; // @[Mux.scala 47:69]
  assign _T_19 = io_expected_out[5] ? 4'h4 : _T_18; // @[Mux.scala 47:69]
  assign _T_20 = io_expected_out[6] ? 4'h3 : _T_19; // @[Mux.scala 47:69]
  assign _T_21 = io_expected_out[7] ? 4'h2 : _T_20; // @[Mux.scala 47:69]
  assign _T_22 = io_expected_out[8] ? 4'h1 : _T_21; // @[Mux.scala 47:69]
  assign _T_23 = io_expected_out[9] ? 4'h0 : _T_22; // @[Mux.scala 47:69]
  assign _GEN_0 = {{15'd0}, io_expected_out[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_24 = _GEN_0 << _T_23; // @[rawFloatFromFN.scala 54:36]
  assign _T_26 = {_T_24[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{2'd0}, _T_23}; // @[rawFloatFromFN.scala 57:26]
  assign _T_27 = _GEN_1 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_28 = _T_3 ? _T_27 : {{1'd0}, io_expected_out[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_29 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{3'd0}, _T_29}; // @[rawFloatFromFN.scala 60:22]
  assign _T_30 = 5'h10 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_30}; // @[rawFloatFromFN.scala 59:15]
  assign _T_32 = _T_28 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_33 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_35 = _T_32[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_38 = _T_35 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_41 = {1'b0,$signed(_T_32)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_43 = _T_3 ? _T_26 : io_expected_out[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_45 = {1'h0,~_T_33,_T_43}; // @[Cat.scala 29:58]
  assign _T_47 = _T_33 ? 3'h0 : _T_41[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_38}; // @[recFNFromFN.scala 48:79]
  assign _T_49 = _T_47 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_52 = {_T_41[2:0],_T_45[9:0]}; // @[Cat.scala 29:58]
  assign _T_53 = {io_expected_out[15],_T_49}; // @[Cat.scala 29:58]
  assign _T_58 = io_actual_out[15:13] == 3'h0; // @[tests.scala 48:26]
  assign _T_60 = io_actual_out[15:13] == 3'h7; // @[tests.scala 48:55]
  assign _T_61 = _T_58 | _T_60; // @[tests.scala 48:39]
  assign _T_62 = io_actual_out[16:13] == io_expected_recOut[16:13]; // @[tests.scala 49:20]
  assign _T_65 = io_actual_out[9:0] == io_expected_recOut[9:0]; // @[tests.scala 49:54]
  assign _T_66 = _T_62 & _T_65; // @[tests.scala 49:31]
  assign _T_68 = io_actual_out[15:13] == 3'h6; // @[tests.scala 50:30]
  assign _T_70 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_71 = _T_68 ? _T_62 : _T_70; // @[tests.scala 50:16]
  assign _T_72 = _T_61 ? _T_66 : _T_71; // @[tests.scala 48:12]
  assign _T_73 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_INToRecFN.scala 80:35]
  assign io_expected_recOut = {_T_53,_T_52}; // @[ValExec_INToRecFN.scala 72:24]
  assign io_actual_out = iNToRecFN_io_out; // @[ValExec_INToRecFN.scala 74:19]
  assign io_actual_exceptionFlags = iNToRecFN_io_exceptionFlags; // @[ValExec_INToRecFN.scala 75:30]
  assign io_check = 1'h1; // @[ValExec_INToRecFN.scala 77:14]
  assign io_pass = _T_72 & _T_73; // @[ValExec_INToRecFN.scala 78:13]
  assign iNToRecFN_io_in = io_in; // @[ValExec_INToRecFN.scala 68:21]
  assign iNToRecFN_io_roundingMode = io_roundingMode; // @[ValExec_INToRecFN.scala 69:33]
endmodule
