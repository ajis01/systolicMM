module MulAddRecFNToRaw_preMul(
  input  [16:0] io_a,
  input  [16:0] io_b,
  input  [16:0] io_c,
  output [10:0] io_mulAddA,
  output [10:0] io_mulAddB,
  output [21:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [6:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [3:0]  io_toPostMul_CDom_CAlignDist,
  output [12:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [11:0] rawA_sig; // @[Cat.scala 29:58]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [11:0] rawB_sig; // @[Cat.scala 29:58]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_36; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire [11:0] rawC_sig; // @[Cat.scala 29:58]
  wire  signProd; // @[MulAddRecFN.scala 98:30]
  wire [7:0] _T_50; // @[MulAddRecFN.scala 101:19]
  wire [7:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  doSubMags; // @[MulAddRecFN.scala 103:30]
  wire [7:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [7:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [6:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _T_57; // @[MulAddRecFN.scala 109:35]
  wire  _T_58; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _T_60; // @[MulAddRecFN.scala 111:60]
  wire  _T_61; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _T_62; // @[MulAddRecFN.scala 115:34]
  wire [5:0] _T_64; // @[MulAddRecFN.scala 115:16]
  wire [5:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [11:0] _T_66; // @[MulAddRecFN.scala 121:16]
  wire [26:0] _T_68; // @[Bitwise.scala 71:12]
  wire [38:0] _T_70; // @[MulAddRecFN.scala 123:11]
  wire [38:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire  _T_74; // @[primitives.scala 121:54]
  wire  _T_76; // @[primitives.scala 121:54]
  wire  _T_78; // @[primitives.scala 124:57]
  wire [2:0] _T_80; // @[primitives.scala 125:20]
  wire [16:0] _T_82; // @[primitives.scala 77:58]
  wire [1:0] _T_86; // @[Cat.scala 29:58]
  wire [2:0] _GEN_1; // @[MulAddRecFN.scala 125:68]
  wire [2:0] _T_87; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _T_90; // @[MulAddRecFN.scala 137:39]
  wire  _T_92; // @[MulAddRecFN.scala 137:44]
  wire  _T_94; // @[MulAddRecFN.scala 138:39]
  wire  _T_95; // @[MulAddRecFN.scala 138:44]
  wire  _T_96; // @[MulAddRecFN.scala 136:16]
  wire [35:0] _T_97; // @[Cat.scala 29:58]
  wire [36:0] alignedSigC; // @[Cat.scala 29:58]
  wire  _T_101; // @[common.scala 81:46]
  wire  _T_104; // @[common.scala 81:46]
  wire  _T_105; // @[MulAddRecFN.scala 149:32]
  wire  _T_108; // @[common.scala 81:46]
  wire [7:0] _T_113; // @[MulAddRecFN.scala 161:53]
  wire [7:0] _T_114; // @[MulAddRecFN.scala 161:12]
  assign rawA_isZero = io_a[15:13] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_4 = io_a[15:14] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA_isNaN = _T_4 & io_a[13]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA_sign = io_a[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA_sExp = {1'b0,$signed(io_a[15:10])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_sig = {1'h0,~rawA_isZero,io_a[9:0]}; // @[Cat.scala 29:58]
  assign rawB_isZero = io_b[15:13] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_20 = io_b[15:14] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB_isNaN = _T_20 & io_b[13]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB_sign = io_b[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB_sExp = {1'b0,$signed(io_b[15:10])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_sig = {1'h0,~rawB_isZero,io_b[9:0]}; // @[Cat.scala 29:58]
  assign rawC_isZero = io_c[15:13] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign _T_36 = io_c[15:14] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC_isNaN = _T_36 & io_c[13]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC_sign = io_c[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC_sExp = {1'b0,$signed(io_c[15:10])}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_sig = {1'h0,~rawC_isZero,io_c[9:0]}; // @[Cat.scala 29:58]
  assign signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  assign _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_T_50) - 8'sh12; // @[MulAddRecFN.scala 101:32]
  assign doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  assign _GEN_0 = {{1{rawC_sExp[6]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[6:0]; // @[MulAddRecFN.scala 108:42]
  assign _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _T_58 = $signed(sNatCAlignDist) < 8'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50]
  assign _T_60 = posNatCAlignDist <= 7'hb; // @[MulAddRecFN.scala 111:60]
  assign _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 111:23]
  assign _T_62 = posNatCAlignDist < 7'h23; // @[MulAddRecFN.scala 115:34]
  assign _T_64 = _T_62 ? posNatCAlignDist[5:0] : 6'h23; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 6'h0 : _T_64; // @[MulAddRecFN.scala 113:12]
  assign _T_66 = doSubMags ? ~rawC_sig : rawC_sig; // @[MulAddRecFN.scala 121:16]
  assign _T_68 = doSubMags ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 71:12]
  assign _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _T_74 = rawC_sig[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_76 = rawC_sig[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_78 = rawC_sig[11:8] != 4'h0; // @[primitives.scala 124:57]
  assign _T_80 = {_T_78,_T_76,_T_74}; // @[primitives.scala 125:20]
  assign _T_82 = -17'sh10000 >>> CAlignDist[5:2]; // @[primitives.scala 77:58]
  assign _T_86 = {_T_82[8],_T_82[9]}; // @[Cat.scala 29:58]
  assign _GEN_1 = {{1'd0}, _T_86}; // @[MulAddRecFN.scala 125:68]
  assign _T_87 = _T_80 & _GEN_1; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = _T_87 != 3'h0; // @[MulAddRecFN.scala 133:11]
  assign _T_90 = mainAlignedSigC[2:0] == 3'h7; // @[MulAddRecFN.scala 137:39]
  assign _T_92 = _T_90 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _T_94 = mainAlignedSigC[2:0] != 3'h0; // @[MulAddRecFN.scala 138:39]
  assign _T_95 = _T_94 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign _T_96 = doSubMags ? _T_92 : _T_95; // @[MulAddRecFN.scala 136:16]
  assign _T_97 = mainAlignedSigC[38:3]; // @[Cat.scala 29:58]
  assign alignedSigC = {_T_97,_T_96}; // @[Cat.scala 29:58]
  assign _T_101 = rawA_isNaN & ~rawA_sig[9]; // @[common.scala 81:46]
  assign _T_104 = rawB_isNaN & ~rawB_sig[9]; // @[common.scala 81:46]
  assign _T_105 = _T_101 | _T_104; // @[MulAddRecFN.scala 149:32]
  assign _T_108 = rawC_isNaN & ~rawC_sig[9]; // @[common.scala 81:46]
  assign _T_113 = $signed(sExpAlignedProd) - 8'shb; // @[MulAddRecFN.scala 161:53]
  assign _T_114 = CIsDominant ? $signed({{1{rawC_sExp[6]}},rawC_sExp}) : $signed(_T_113); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[10:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[10:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[22:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_105 | _T_108; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_4 & ~io_a[13]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[15:13] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_20 & ~io_b[13]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[15:13] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_36 & io_c[13]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_36 & ~io_c[13]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[15:13] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_114[6:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = ~rawC_isZero & _T_61; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[3:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[35:23]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [6:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [3:0]  io_fromPreMul_CDom_CAlignDist,
  input  [12:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [22:0] io_mulAddResult,
  input  [2:0]  io_roundingMode,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [6:0]  io_rawOut_sExp,
  output [13:0] io_rawOut_sig
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [12:0] _T_2; // @[MulAddRecFN.scala 195:47]
  wire [12:0] _T_3; // @[MulAddRecFN.scala 194:16]
  wire [35:0] sigSum; // @[Cat.scala 29:58]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69]
  wire [6:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [6:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [23:0] _T_14; // @[Cat.scala 29:58]
  wire [23:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _T_17; // @[MulAddRecFN.scala 217:36]
  wire  _T_19; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [38:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [38:0] _T_20; // @[MulAddRecFN.scala 221:24]
  wire [15:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire  _T_25; // @[primitives.scala 121:54]
  wire  _T_27; // @[primitives.scala 121:54]
  wire  _T_29; // @[primitives.scala 124:57]
  wire [2:0] _T_31; // @[primitives.scala 125:20]
  wire [4:0] _T_34; // @[primitives.scala 77:58]
  wire [1:0] _T_38; // @[Cat.scala 29:58]
  wire [2:0] _GEN_2; // @[MulAddRecFN.scala 224:72]
  wire [2:0] _T_39; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire  _T_42; // @[MulAddRecFN.scala 228:32]
  wire  _T_43; // @[MulAddRecFN.scala 228:36]
  wire  _T_44; // @[MulAddRecFN.scala 228:61]
  wire [13:0] CDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [24:0] _GEN_3; // @[MulAddRecFN.scala 238:41]
  wire [24:0] _T_49; // @[MulAddRecFN.scala 238:41]
  wire [24:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  _T_52; // @[primitives.scala 104:54]
  wire  _T_54; // @[primitives.scala 104:54]
  wire  _T_56; // @[primitives.scala 104:54]
  wire  _T_58; // @[primitives.scala 104:54]
  wire  _T_60; // @[primitives.scala 104:54]
  wire  _T_62; // @[primitives.scala 104:54]
  wire  _T_64; // @[primitives.scala 104:54]
  wire  _T_66; // @[primitives.scala 104:54]
  wire  _T_68; // @[primitives.scala 104:54]
  wire  _T_70; // @[primitives.scala 104:54]
  wire  _T_72; // @[primitives.scala 104:54]
  wire  _T_74; // @[primitives.scala 104:54]
  wire [5:0] _T_81; // @[primitives.scala 108:20]
  wire [12:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [3:0] _T_101; // @[Mux.scala 47:69]
  wire [3:0] _T_102; // @[Mux.scala 47:69]
  wire [3:0] _T_103; // @[Mux.scala 47:69]
  wire [3:0] _T_104; // @[Mux.scala 47:69]
  wire [3:0] _T_105; // @[Mux.scala 47:69]
  wire [3:0] _T_106; // @[Mux.scala 47:69]
  wire [3:0] _T_107; // @[Mux.scala 47:69]
  wire [3:0] _T_108; // @[Mux.scala 47:69]
  wire [3:0] _T_109; // @[Mux.scala 47:69]
  wire [3:0] _T_110; // @[Mux.scala 47:69]
  wire [3:0] _T_111; // @[Mux.scala 47:69]
  wire [3:0] notCDom_normDistReduced2; // @[Mux.scala 47:69]
  wire [4:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [5:0] _T_112; // @[MulAddRecFN.scala 243:69]
  wire [6:0] _GEN_4; // @[MulAddRecFN.scala 243:46]
  wire [6:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [55:0] _GEN_5; // @[MulAddRecFN.scala 245:27]
  wire [55:0] _T_115; // @[MulAddRecFN.scala 245:27]
  wire [15:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire [6:0] _T_117; // @[MulAddRecFN.scala 249:55]
  wire  _T_120; // @[primitives.scala 104:54]
  wire  _T_122; // @[primitives.scala 104:54]
  wire  _T_124; // @[primitives.scala 104:54]
  wire [3:0] _T_129; // @[primitives.scala 108:20]
  wire [8:0] _T_132; // @[primitives.scala 77:58]
  wire [2:0] _T_139; // @[Cat.scala 29:58]
  wire [3:0] _GEN_6; // @[MulAddRecFN.scala 249:78]
  wire [3:0] _T_140; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire  _T_143; // @[MulAddRecFN.scala 254:35]
  wire  _T_144; // @[MulAddRecFN.scala 254:39]
  wire [13:0] notCDom_sig; // @[Cat.scala 29:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _T_146; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _T_147; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _T_148; // @[MulAddRecFN.scala 274:31]
  wire  _T_149; // @[MulAddRecFN.scala 273:35]
  wire  _T_150; // @[MulAddRecFN.scala 275:32]
  wire  _T_151; // @[MulAddRecFN.scala 274:57]
  wire  _T_154; // @[MulAddRecFN.scala 276:36]
  wire  _T_155; // @[MulAddRecFN.scala 277:61]
  wire  _T_156; // @[MulAddRecFN.scala 278:35]
  wire  _T_160; // @[MulAddRecFN.scala 285:42]
  wire  _T_162; // @[MulAddRecFN.scala 287:27]
  wire  _T_163; // @[MulAddRecFN.scala 288:31]
  wire  _T_164; // @[MulAddRecFN.scala 287:54]
  wire  _T_166; // @[MulAddRecFN.scala 289:26]
  wire  _T_167; // @[MulAddRecFN.scala 289:48]
  wire  _T_168; // @[MulAddRecFN.scala 290:36]
  wire  _T_169; // @[MulAddRecFN.scala 288:43]
  wire  _T_170; // @[MulAddRecFN.scala 291:26]
  wire  _T_171; // @[MulAddRecFN.scala 292:37]
  wire  _T_172; // @[MulAddRecFN.scala 291:46]
  wire  _T_173; // @[MulAddRecFN.scala 290:48]
  wire  _T_176; // @[MulAddRecFN.scala 293:28]
  wire  _T_177; // @[MulAddRecFN.scala 294:17]
  wire  _T_178; // @[MulAddRecFN.scala 293:49]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 13'h1; // @[MulAddRecFN.scala 195:47]
  assign _T_3 = io_mulAddResult[22] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum = {_T_3,io_mulAddResult[21:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{5{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[12:11],sigSum[33:13]}; // @[Cat.scala 29:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[35:12] : _T_14; // @[MulAddRecFN.scala 207:12]
  assign _T_17 = ~sigSum[11:1] != 11'h0; // @[MulAddRecFN.scala 217:36]
  assign _T_19 = sigSum[12:1] != 12'h0; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{15'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _T_20[23:8]; // @[MulAddRecFN.scala 221:56]
  assign _T_25 = CDom_absSigSum[3:0] != 4'h0; // @[primitives.scala 121:54]
  assign _T_27 = CDom_absSigSum[7:4] != 4'h0; // @[primitives.scala 121:54]
  assign _T_29 = CDom_absSigSum[10:8] != 3'h0; // @[primitives.scala 124:57]
  assign _T_31 = {_T_29,_T_27,_T_25}; // @[primitives.scala 125:20]
  assign _T_34 = -5'sh10 >>> ~io_fromPreMul_CDom_CAlignDist[3:2]; // @[primitives.scala 77:58]
  assign _T_38 = {_T_34[1],_T_34[2]}; // @[Cat.scala 29:58]
  assign _GEN_2 = {{1'd0}, _T_38}; // @[MulAddRecFN.scala 224:72]
  assign _T_39 = _T_31 & _GEN_2; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = _T_39 != 3'h0; // @[MulAddRecFN.scala 225:73]
  assign _T_42 = CDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 228:32]
  assign _T_43 = _T_42 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign _T_44 = _T_43 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_mainSig[15:3],_T_44}; // @[Cat.scala 29:58]
  assign notCDom_signSigSum = sigSum[25]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_3 = {{24'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _T_49 = sigSum[24:0] + _GEN_3; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[24:0] : _T_49; // @[MulAddRecFN.scala 236:12]
  assign _T_52 = notCDom_absSigSum[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_54 = notCDom_absSigSum[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_56 = notCDom_absSigSum[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_58 = notCDom_absSigSum[7:6] != 2'h0; // @[primitives.scala 104:54]
  assign _T_60 = notCDom_absSigSum[9:8] != 2'h0; // @[primitives.scala 104:54]
  assign _T_62 = notCDom_absSigSum[11:10] != 2'h0; // @[primitives.scala 104:54]
  assign _T_64 = notCDom_absSigSum[13:12] != 2'h0; // @[primitives.scala 104:54]
  assign _T_66 = notCDom_absSigSum[15:14] != 2'h0; // @[primitives.scala 104:54]
  assign _T_68 = notCDom_absSigSum[17:16] != 2'h0; // @[primitives.scala 104:54]
  assign _T_70 = notCDom_absSigSum[19:18] != 2'h0; // @[primitives.scala 104:54]
  assign _T_72 = notCDom_absSigSum[21:20] != 2'h0; // @[primitives.scala 104:54]
  assign _T_74 = notCDom_absSigSum[23:22] != 2'h0; // @[primitives.scala 104:54]
  assign _T_81 = {_T_62,_T_60,_T_58,_T_56,_T_54,_T_52}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {notCDom_absSigSum[24],_T_74,_T_72,_T_70,_T_68,_T_66,_T_64,_T_81}; // @[primitives.scala 108:20]
  assign _T_101 = notCDom_reduced2AbsSigSum[1] ? 4'hb : 4'hc; // @[Mux.scala 47:69]
  assign _T_102 = notCDom_reduced2AbsSigSum[2] ? 4'ha : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = notCDom_reduced2AbsSigSum[3] ? 4'h9 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = notCDom_reduced2AbsSigSum[4] ? 4'h8 : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = notCDom_reduced2AbsSigSum[5] ? 4'h7 : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = notCDom_reduced2AbsSigSum[6] ? 4'h6 : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = notCDom_reduced2AbsSigSum[7] ? 4'h5 : _T_106; // @[Mux.scala 47:69]
  assign _T_108 = notCDom_reduced2AbsSigSum[8] ? 4'h4 : _T_107; // @[Mux.scala 47:69]
  assign _T_109 = notCDom_reduced2AbsSigSum[9] ? 4'h3 : _T_108; // @[Mux.scala 47:69]
  assign _T_110 = notCDom_reduced2AbsSigSum[10] ? 4'h2 : _T_109; // @[Mux.scala 47:69]
  assign _T_111 = notCDom_reduced2AbsSigSum[11] ? 4'h1 : _T_110; // @[Mux.scala 47:69]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[12] ? 4'h0 : _T_111; // @[Mux.scala 47:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _T_112 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_4 = {{1{_T_112[5]}},_T_112}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46]
  assign _GEN_5 = {{31'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _T_115 = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _T_115[25:10]; // @[MulAddRecFN.scala 245:50]
  assign _T_117 = {notCDom_reduced2AbsSigSum[5:0], 1'h0}; // @[MulAddRecFN.scala 249:55]
  assign _T_120 = _T_117[1:0] != 2'h0; // @[primitives.scala 104:54]
  assign _T_122 = _T_117[3:2] != 2'h0; // @[primitives.scala 104:54]
  assign _T_124 = _T_117[5:4] != 2'h0; // @[primitives.scala 104:54]
  assign _T_129 = {_T_117[6],_T_124,_T_122,_T_120}; // @[primitives.scala 108:20]
  assign _T_132 = -9'sh100 >>> ~notCDom_normDistReduced2[3:1]; // @[primitives.scala 77:58]
  assign _T_139 = {_T_132[1],_T_132[2],_T_132[3]}; // @[Cat.scala 29:58]
  assign _GEN_6 = {{1'd0}, _T_139}; // @[MulAddRecFN.scala 249:78]
  assign _T_140 = _T_129 & _GEN_6; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = _T_140 != 4'h0; // @[MulAddRecFN.scala 251:11]
  assign _T_143 = notCDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 254:35]
  assign _T_144 = _T_143 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_mainSig[15:3],_T_144}; // @[Cat.scala 29:58]
  assign notCDom_completeCancellation = notCDom_sig[13:12] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _T_146 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_146; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _T_147 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _T_147 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _T_148 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _T_149 = io_fromPreMul_isSigNaNAny | _T_148; // @[MulAddRecFN.scala 273:35]
  assign _T_150 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _T_151 = _T_149 | _T_150; // @[MulAddRecFN.scala 274:57]
  assign _T_154 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _T_155 = _T_154 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _T_156 = _T_155 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _T_160 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _T_162 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _T_163 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _T_164 = _T_162 | _T_163; // @[MulAddRecFN.scala 287:54]
  assign _T_166 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _T_167 = _T_166 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _T_168 = _T_167 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _T_169 = _T_164 | _T_168; // @[MulAddRecFN.scala 288:43]
  assign _T_170 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _T_171 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _T_172 = _T_170 & _T_171; // @[MulAddRecFN.scala 291:46]
  assign _T_173 = _T_169 | _T_172; // @[MulAddRecFN.scala 290:48]
  assign _T_176 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _T_177 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _T_178 = _T_176 & _T_177; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_151 | _T_156; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_160; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_173 | _T_178; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [6:0]  io_in_sExp,
  input  [13:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [16:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire [64:0] _T_5; // @[primitives.scala 77:58]
  wire [7:0] _T_11; // @[Bitwise.scala 102:31]
  wire [7:0] _T_13; // @[Bitwise.scala 102:65]
  wire [7:0] _T_15; // @[Bitwise.scala 102:75]
  wire [7:0] _T_16; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_0; // @[Bitwise.scala 102:31]
  wire [7:0] _T_21; // @[Bitwise.scala 102:31]
  wire [7:0] _T_23; // @[Bitwise.scala 102:65]
  wire [7:0] _T_25; // @[Bitwise.scala 102:75]
  wire [7:0] _T_26; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [7:0] _T_31; // @[Bitwise.scala 102:31]
  wire [7:0] _T_33; // @[Bitwise.scala 102:65]
  wire [7:0] _T_35; // @[Bitwise.scala 102:75]
  wire [7:0] _T_36; // @[Bitwise.scala 102:39]
  wire [11:0] _T_47; // @[Cat.scala 29:58]
  wire [11:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [11:0] _T_48; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [13:0] _T_49; // @[Cat.scala 29:58]
  wire [13:0] _T_51; // @[Cat.scala 29:58]
  wire [13:0] _T_53; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [13:0] _T_54; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_55; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [13:0] _T_56; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_57; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_58; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _T_59; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _T_60; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _T_61; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  _T_62; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [13:0] _T_63; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [12:0] _T_65; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _T_66; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _T_68; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [12:0] _T_70; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [12:0] _T_72; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [13:0] _T_74; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _T_76; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [12:0] _T_78; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [12:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] _T_79; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] _T_80; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _T_82; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [6:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [7:0] _T_83; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [5:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [9:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_88; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  _T_93; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _T_95; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _T_97; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _T_98; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _T_100; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _T_101; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  _T_102; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  _T_105; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _T_106; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _T_107; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _T_108; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _T_111; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _T_112; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _T_116; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _T_118; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _T_119; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _T_120; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _T_121; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _T_123; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _T_128; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _T_130; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _T_132; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _T_133; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _T_135; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_136; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [5:0] _T_137; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [5:0] _T_139; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [5:0] _T_141; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [5:0] _T_143; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [5:0] _T_144; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [5:0] _T_146; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [5:0] _T_147; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [5:0] _T_149; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [5:0] _T_150; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [5:0] _T_151; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [5:0] _T_152; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [5:0] _T_153; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [5:0] _T_154; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [5:0] _T_155; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [5:0] _T_156; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [5:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_157; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_158; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [9:0] _T_159; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [9:0] _T_160; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] _T_162; // @[Bitwise.scala 71:12]
  wire [9:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [6:0] _T_163; // @[Cat.scala 29:58]
  wire [1:0] _T_165; // @[Cat.scala 29:58]
  wire [2:0] _T_167; // @[Cat.scala 29:58]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[13]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign _T_5 = -65'sh10000000000000000 >>> ~io_in_sExp[5:0]; // @[primitives.scala 77:58]
  assign _T_11 = {{4'd0}, _T_5[14:11]}; // @[Bitwise.scala 102:31]
  assign _T_13 = {_T_5[10:7], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_15 = _T_13 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_16 = _T_11 | _T_15; // @[Bitwise.scala 102:39]
  assign _GEN_0 = {{2'd0}, _T_16[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_21 = _GEN_0 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_23 = {_T_16[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_25 = _T_23 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_26 = _T_21 | _T_25; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{1'd0}, _T_26[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_31 = _GEN_1 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_33 = {_T_26[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_35 = _T_33 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_36 = _T_31 | _T_35; // @[Bitwise.scala 102:39]
  assign _T_47 = {_T_36,_T_5[15],_T_5[16],_T_5[17],_T_5[18]}; // @[Cat.scala 29:58]
  assign _GEN_2 = {{11'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_48 = _T_47 | _GEN_2; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign _T_49 = {_T_48,2'h3}; // @[Cat.scala 29:58]
  assign _T_51 = {1'h0,_T_49[13:1]}; // @[Cat.scala 29:58]
  assign _T_53 = ~_T_51 & _T_49; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _T_54 = io_in_sig & _T_53; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign _T_55 = _T_54 != 14'h0; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _T_56 = io_in_sig & _T_51; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign _T_57 = _T_56 != 14'h0; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign _T_58 = _T_55 | _T_57; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _T_59 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _T_60 = _T_59 & _T_55; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _T_61 = roundMagUp & _T_58; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign _T_62 = _T_60 | _T_61; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _T_63 = io_in_sig | _T_49; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _T_65 = _T_63[13:2] + 12'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _T_66 = roundingMode_near_even & _T_55; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _T_68 = _T_66 & ~_T_57; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _T_70 = _T_68 ? _T_49[13:1] : 13'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _T_72 = _T_65 & ~_T_70; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _T_74 = io_in_sig & ~_T_49; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _T_76 = roundingMode_odd & _T_58; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _T_78 = _T_76 ? _T_53[13:1] : 13'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_3 = {{1'd0}, _T_74[13:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_79 = _GEN_3 | _T_78; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _T_80 = _T_62 ? _T_72 : _T_79; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _T_82 = {1'b0,$signed(_T_80[12:11])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_4 = {{4{_T_82[2]}},_T_82}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign _T_83 = $signed(io_in_sExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = _T_83[5:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? _T_80[10:1] : _T_80[9:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _T_88 = _T_83[7:4]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_T_88) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(_T_83) < 8'sh8; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign _T_93 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _T_95 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _T_97 = io_in_sig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _T_98 = _T_95 | _T_97; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _T_100 = _T_59 & _T_93; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _T_101 = roundMagUp & _T_98; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign _T_102 = _T_100 | _T_101; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign _T_105 = doShiftSigDown1 ? _T_80[12] : _T_80[11]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _T_106 = io_in_sExp[6:5]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _T_107 = $signed(_T_106) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _T_108 = _T_58 & _T_107; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _T_111 = doShiftSigDown1 ? _T_49[3] : _T_49[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _T_112 = _T_108 & _T_111; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _T_116 = doShiftSigDown1 ? _T_49[4] : _T_49[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _T_118 = io_detectTininess & ~_T_116; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _T_119 = _T_118 & _T_105; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _T_120 = _T_119 & _T_55; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _T_121 = _T_120 & _T_102; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _T_123 = _T_112 & ~_T_121; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _T_123; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | _T_58; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign _T_128 = ~isNaNOut & ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _T_128 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _T_130 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _T_130; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _T_59 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _T_132 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _T_133 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _T_132 & _T_133; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _T_135 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = io_in_isInf | _T_135; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _T_136 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _T_137 = _T_136 ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _T_139 = common_expOut & ~_T_137; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _T_141 = pegMinNonzeroMagOut ? 6'h37 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _T_143 = _T_139 & ~_T_141; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _T_144 = pegMaxFiniteMagOut ? 6'h10 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _T_146 = _T_143 & ~_T_144; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _T_147 = notNaN_isInfOut ? 6'h8 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _T_149 = _T_146 & ~_T_147; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _T_150 = pegMinNonzeroMagOut ? 6'h8 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _T_151 = _T_149 | _T_150; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _T_152 = pegMaxFiniteMagOut ? 6'h2f : 6'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _T_153 = _T_151 | _T_152; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _T_154 = notNaN_isInfOut ? 6'h30 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _T_155 = _T_153 | _T_154; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _T_156 = isNaNOut ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _T_155 | _T_156; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _T_157 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _T_158 = _T_157 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _T_159 = isNaNOut ? 10'h200 : 10'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _T_160 = _T_158 ? _T_159 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_162 = pegMaxFiniteMagOut ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign fractOut = _T_160 | _T_162; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign _T_163 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign _T_165 = {underflow,inexact}; // @[Cat.scala 29:58]
  assign _T_167 = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 29:58]
  assign io_out = {_T_163,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {_T_167,_T_165}; // @[RoundAnyRawFNToRecFN.scala 285:23]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [6:0]  io_in_sExp,
  input  [13:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [16:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [6:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [13:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [16:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
endmodule
module MulAddRecFN(
  input  [16:0] io_a,
  input  [16:0] io_b,
  input  [16:0] io_c,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [16:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire [16:0] mulAddRecFNToRaw_preMul_io_a; // @[MulAddRecFN.scala 318:15]
  wire [16:0] mulAddRecFNToRaw_preMul_io_b; // @[MulAddRecFN.scala 318:15]
  wire [16:0] mulAddRecFNToRaw_preMul_io_c; // @[MulAddRecFN.scala 318:15]
  wire [10:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[MulAddRecFN.scala 318:15]
  wire [10:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 318:15]
  wire [21:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 318:15]
  wire [6:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 318:15]
  wire [3:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 318:15]
  wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 320:15]
  wire [6:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 320:15]
  wire [3:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 320:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire [22:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[MulAddRecFN.scala 320:15]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 320:15]
  wire [6:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 320:15]
  wire [13:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 320:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulAddRecFN.scala 340:15]
  wire [6:0] roundRawFNToRecFN_io_in_sExp; // @[MulAddRecFN.scala 340:15]
  wire [13:0] roundRawFNToRecFN_io_in_sig; // @[MulAddRecFN.scala 340:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[MulAddRecFN.scala 340:15]
  wire [16:0] roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 340:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[MulAddRecFN.scala 340:15]
  wire [21:0] _T; // @[MulAddRecFN.scala 328:45]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[MulAddRecFN.scala 318:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[MulAddRecFN.scala 320:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[MulAddRecFN.scala 340:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags)
  );
  assign _T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 328:45]
  assign io_out = roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 346:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[MulAddRecFN.scala 347:23]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[MulAddRecFN.scala 323:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[MulAddRecFN.scala 324:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[MulAddRecFN.scala 325:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 334:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = io_roundingMode; // @[MulAddRecFN.scala 335:46]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 341:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_roundingMode = io_roundingMode; // @[MulAddRecFN.scala 344:39]
  assign roundRawFNToRecFN_io_detectTininess = io_detectTininess; // @[MulAddRecFN.scala 345:41]
endmodule
module ValExec_MulAddRecF16(
  input         clock,
  input         reset,
  input  [15:0] io_a,
  input  [15:0] io_b,
  input  [15:0] io_c,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [15:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [16:0] io_expected_recOut,
  output [16:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [16:0] mulAddRecFN_io_a; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [16:0] mulAddRecFN_io_b; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [16:0] mulAddRecFN_io_c; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [2:0] mulAddRecFN_io_roundingMode; // @[ValExec_MulAddRecFN.scala 66:29]
  wire  mulAddRecFN_io_detectTininess; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [16:0] mulAddRecFN_io_out; // @[ValExec_MulAddRecFN.scala 66:29]
  wire [4:0] mulAddRecFN_io_exceptionFlags; // @[ValExec_MulAddRecFN.scala 66:29]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_15; // @[Mux.scala 47:69]
  wire [3:0] _T_16; // @[Mux.scala 47:69]
  wire [3:0] _T_17; // @[Mux.scala 47:69]
  wire [3:0] _T_18; // @[Mux.scala 47:69]
  wire [3:0] _T_19; // @[Mux.scala 47:69]
  wire [3:0] _T_20; // @[Mux.scala 47:69]
  wire [3:0] _T_21; // @[Mux.scala 47:69]
  wire [3:0] _T_22; // @[Mux.scala 47:69]
  wire [3:0] _T_23; // @[Mux.scala 47:69]
  wire [24:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_24; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_26; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_27; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_28; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_29; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_30; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_32; // @[rawFloatFromFN.scala 59:15]
  wire  _T_33; // @[rawFloatFromFN.scala 62:34]
  wire  _T_35; // @[rawFloatFromFN.scala 63:62]
  wire  _T_38; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_41; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_43; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_45; // @[Cat.scala 29:58]
  wire [2:0] _T_47; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_49; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_52; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[Cat.scala 29:58]
  wire  _T_58; // @[rawFloatFromFN.scala 50:34]
  wire  _T_59; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_70; // @[Mux.scala 47:69]
  wire [3:0] _T_71; // @[Mux.scala 47:69]
  wire [3:0] _T_72; // @[Mux.scala 47:69]
  wire [3:0] _T_73; // @[Mux.scala 47:69]
  wire [3:0] _T_74; // @[Mux.scala 47:69]
  wire [3:0] _T_75; // @[Mux.scala 47:69]
  wire [3:0] _T_76; // @[Mux.scala 47:69]
  wire [3:0] _T_77; // @[Mux.scala 47:69]
  wire [3:0] _T_78; // @[Mux.scala 47:69]
  wire [24:0] _GEN_5; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_79; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_81; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_6; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_82; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_83; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_84; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_85; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_87; // @[rawFloatFromFN.scala 59:15]
  wire  _T_88; // @[rawFloatFromFN.scala 62:34]
  wire  _T_90; // @[rawFloatFromFN.scala 63:62]
  wire  _T_93; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_96; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_98; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_100; // @[Cat.scala 29:58]
  wire [2:0] _T_102; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_104; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_107; // @[Cat.scala 29:58]
  wire [3:0] _T_108; // @[Cat.scala 29:58]
  wire  _T_113; // @[rawFloatFromFN.scala 50:34]
  wire  _T_114; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_125; // @[Mux.scala 47:69]
  wire [3:0] _T_126; // @[Mux.scala 47:69]
  wire [3:0] _T_127; // @[Mux.scala 47:69]
  wire [3:0] _T_128; // @[Mux.scala 47:69]
  wire [3:0] _T_129; // @[Mux.scala 47:69]
  wire [3:0] _T_130; // @[Mux.scala 47:69]
  wire [3:0] _T_131; // @[Mux.scala 47:69]
  wire [3:0] _T_132; // @[Mux.scala 47:69]
  wire [3:0] _T_133; // @[Mux.scala 47:69]
  wire [24:0] _GEN_10; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_134; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_136; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_11; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_137; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_138; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_139; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_12; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_140; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_13; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_142; // @[rawFloatFromFN.scala 59:15]
  wire  _T_143; // @[rawFloatFromFN.scala 62:34]
  wire  _T_145; // @[rawFloatFromFN.scala 63:62]
  wire  _T_148; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_151; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_153; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_155; // @[Cat.scala 29:58]
  wire [2:0] _T_157; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_14; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_159; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_162; // @[Cat.scala 29:58]
  wire [3:0] _T_163; // @[Cat.scala 29:58]
  wire  _T_168; // @[rawFloatFromFN.scala 50:34]
  wire  _T_169; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _T_180; // @[Mux.scala 47:69]
  wire [3:0] _T_181; // @[Mux.scala 47:69]
  wire [3:0] _T_182; // @[Mux.scala 47:69]
  wire [3:0] _T_183; // @[Mux.scala 47:69]
  wire [3:0] _T_184; // @[Mux.scala 47:69]
  wire [3:0] _T_185; // @[Mux.scala 47:69]
  wire [3:0] _T_186; // @[Mux.scala 47:69]
  wire [3:0] _T_187; // @[Mux.scala 47:69]
  wire [3:0] _T_188; // @[Mux.scala 47:69]
  wire [24:0] _GEN_15; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _T_189; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] _T_191; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_16; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_192; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _T_193; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_194; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_17; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _T_195; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_18; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] _T_197; // @[rawFloatFromFN.scala 59:15]
  wire  _T_198; // @[rawFloatFromFN.scala 62:34]
  wire  _T_200; // @[rawFloatFromFN.scala 63:62]
  wire  _T_203; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] _T_206; // @[rawFloatFromFN.scala 70:48]
  wire [9:0] _T_208; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] _T_210; // @[Cat.scala 29:58]
  wire [2:0] _T_212; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_19; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_214; // @[recFNFromFN.scala 48:79]
  wire [12:0] _T_217; // @[Cat.scala 29:58]
  wire [3:0] _T_218; // @[Cat.scala 29:58]
  wire  _T_223; // @[tests.scala 48:26]
  wire  _T_225; // @[tests.scala 48:55]
  wire  _T_226; // @[tests.scala 48:39]
  wire  _T_227; // @[tests.scala 49:20]
  wire  _T_230; // @[tests.scala 49:54]
  wire  _T_231; // @[tests.scala 49:31]
  wire  _T_233; // @[tests.scala 50:30]
  wire  _T_235; // @[tests.scala 50:66]
  wire  _T_236; // @[tests.scala 50:16]
  wire  _T_237; // @[tests.scala 48:12]
  wire  _T_238; // @[ValExec_MulAddRecFN.scala 82:35]
  MulAddRecFN mulAddRecFN ( // @[ValExec_MulAddRecFN.scala 66:29]
    .io_a(mulAddRecFN_io_a),
    .io_b(mulAddRecFN_io_b),
    .io_c(mulAddRecFN_io_c),
    .io_roundingMode(mulAddRecFN_io_roundingMode),
    .io_detectTininess(mulAddRecFN_io_detectTininess),
    .io_out(mulAddRecFN_io_out),
    .io_exceptionFlags(mulAddRecFN_io_exceptionFlags)
  );
  assign _T_3 = io_a[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_a[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_15 = io_a[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_16 = io_a[2] ? 4'h7 : _T_15; // @[Mux.scala 47:69]
  assign _T_17 = io_a[3] ? 4'h6 : _T_16; // @[Mux.scala 47:69]
  assign _T_18 = io_a[4] ? 4'h5 : _T_17; // @[Mux.scala 47:69]
  assign _T_19 = io_a[5] ? 4'h4 : _T_18; // @[Mux.scala 47:69]
  assign _T_20 = io_a[6] ? 4'h3 : _T_19; // @[Mux.scala 47:69]
  assign _T_21 = io_a[7] ? 4'h2 : _T_20; // @[Mux.scala 47:69]
  assign _T_22 = io_a[8] ? 4'h1 : _T_21; // @[Mux.scala 47:69]
  assign _T_23 = io_a[9] ? 4'h0 : _T_22; // @[Mux.scala 47:69]
  assign _GEN_0 = {{15'd0}, io_a[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_24 = _GEN_0 << _T_23; // @[rawFloatFromFN.scala 54:36]
  assign _T_26 = {_T_24[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{2'd0}, _T_23}; // @[rawFloatFromFN.scala 57:26]
  assign _T_27 = _GEN_1 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_28 = _T_3 ? _T_27 : {{1'd0}, io_a[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_29 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{3'd0}, _T_29}; // @[rawFloatFromFN.scala 60:22]
  assign _T_30 = 5'h10 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_30}; // @[rawFloatFromFN.scala 59:15]
  assign _T_32 = _T_28 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_33 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_35 = _T_32[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_38 = _T_35 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_41 = {1'b0,$signed(_T_32)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_43 = _T_3 ? _T_26 : io_a[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_45 = {1'h0,~_T_33,_T_43}; // @[Cat.scala 29:58]
  assign _T_47 = _T_33 ? 3'h0 : _T_41[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_38}; // @[recFNFromFN.scala 48:79]
  assign _T_49 = _T_47 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_52 = {_T_41[2:0],_T_45[9:0]}; // @[Cat.scala 29:58]
  assign _T_53 = {io_a[15],_T_49}; // @[Cat.scala 29:58]
  assign _T_58 = io_b[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_59 = io_b[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_70 = io_b[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_71 = io_b[2] ? 4'h7 : _T_70; // @[Mux.scala 47:69]
  assign _T_72 = io_b[3] ? 4'h6 : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = io_b[4] ? 4'h5 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = io_b[5] ? 4'h4 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = io_b[6] ? 4'h3 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = io_b[7] ? 4'h2 : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = io_b[8] ? 4'h1 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = io_b[9] ? 4'h0 : _T_77; // @[Mux.scala 47:69]
  assign _GEN_5 = {{15'd0}, io_b[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_79 = _GEN_5 << _T_78; // @[rawFloatFromFN.scala 54:36]
  assign _T_81 = {_T_79[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_6 = {{2'd0}, _T_78}; // @[rawFloatFromFN.scala 57:26]
  assign _T_82 = _GEN_6 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_83 = _T_58 ? _T_82 : {{1'd0}, io_b[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_84 = _T_58 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_7 = {{3'd0}, _T_84}; // @[rawFloatFromFN.scala 60:22]
  assign _T_85 = 5'h10 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_8 = {{1'd0}, _T_85}; // @[rawFloatFromFN.scala 59:15]
  assign _T_87 = _T_83 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  assign _T_88 = _T_58 & _T_59; // @[rawFloatFromFN.scala 62:34]
  assign _T_90 = _T_87[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_93 = _T_90 & ~_T_59; // @[rawFloatFromFN.scala 66:33]
  assign _T_96 = {1'b0,$signed(_T_87)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_98 = _T_58 ? _T_81 : io_b[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_100 = {1'h0,~_T_88,_T_98}; // @[Cat.scala 29:58]
  assign _T_102 = _T_88 ? 3'h0 : _T_96[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_9 = {{2'd0}, _T_93}; // @[recFNFromFN.scala 48:79]
  assign _T_104 = _T_102 | _GEN_9; // @[recFNFromFN.scala 48:79]
  assign _T_107 = {_T_96[2:0],_T_100[9:0]}; // @[Cat.scala 29:58]
  assign _T_108 = {io_b[15],_T_104}; // @[Cat.scala 29:58]
  assign _T_113 = io_c[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_114 = io_c[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_125 = io_c[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_126 = io_c[2] ? 4'h7 : _T_125; // @[Mux.scala 47:69]
  assign _T_127 = io_c[3] ? 4'h6 : _T_126; // @[Mux.scala 47:69]
  assign _T_128 = io_c[4] ? 4'h5 : _T_127; // @[Mux.scala 47:69]
  assign _T_129 = io_c[5] ? 4'h4 : _T_128; // @[Mux.scala 47:69]
  assign _T_130 = io_c[6] ? 4'h3 : _T_129; // @[Mux.scala 47:69]
  assign _T_131 = io_c[7] ? 4'h2 : _T_130; // @[Mux.scala 47:69]
  assign _T_132 = io_c[8] ? 4'h1 : _T_131; // @[Mux.scala 47:69]
  assign _T_133 = io_c[9] ? 4'h0 : _T_132; // @[Mux.scala 47:69]
  assign _GEN_10 = {{15'd0}, io_c[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_134 = _GEN_10 << _T_133; // @[rawFloatFromFN.scala 54:36]
  assign _T_136 = {_T_134[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_11 = {{2'd0}, _T_133}; // @[rawFloatFromFN.scala 57:26]
  assign _T_137 = _GEN_11 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_138 = _T_113 ? _T_137 : {{1'd0}, io_c[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_139 = _T_113 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_12 = {{3'd0}, _T_139}; // @[rawFloatFromFN.scala 60:22]
  assign _T_140 = 5'h10 | _GEN_12; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_13 = {{1'd0}, _T_140}; // @[rawFloatFromFN.scala 59:15]
  assign _T_142 = _T_138 + _GEN_13; // @[rawFloatFromFN.scala 59:15]
  assign _T_143 = _T_113 & _T_114; // @[rawFloatFromFN.scala 62:34]
  assign _T_145 = _T_142[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_148 = _T_145 & ~_T_114; // @[rawFloatFromFN.scala 66:33]
  assign _T_151 = {1'b0,$signed(_T_142)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_153 = _T_113 ? _T_136 : io_c[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_155 = {1'h0,~_T_143,_T_153}; // @[Cat.scala 29:58]
  assign _T_157 = _T_143 ? 3'h0 : _T_151[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_14 = {{2'd0}, _T_148}; // @[recFNFromFN.scala 48:79]
  assign _T_159 = _T_157 | _GEN_14; // @[recFNFromFN.scala 48:79]
  assign _T_162 = {_T_151[2:0],_T_155[9:0]}; // @[Cat.scala 29:58]
  assign _T_163 = {io_c[15],_T_159}; // @[Cat.scala 29:58]
  assign _T_168 = io_expected_out[14:10] == 5'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_169 = io_expected_out[9:0] == 10'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_180 = io_expected_out[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  assign _T_181 = io_expected_out[2] ? 4'h7 : _T_180; // @[Mux.scala 47:69]
  assign _T_182 = io_expected_out[3] ? 4'h6 : _T_181; // @[Mux.scala 47:69]
  assign _T_183 = io_expected_out[4] ? 4'h5 : _T_182; // @[Mux.scala 47:69]
  assign _T_184 = io_expected_out[5] ? 4'h4 : _T_183; // @[Mux.scala 47:69]
  assign _T_185 = io_expected_out[6] ? 4'h3 : _T_184; // @[Mux.scala 47:69]
  assign _T_186 = io_expected_out[7] ? 4'h2 : _T_185; // @[Mux.scala 47:69]
  assign _T_187 = io_expected_out[8] ? 4'h1 : _T_186; // @[Mux.scala 47:69]
  assign _T_188 = io_expected_out[9] ? 4'h0 : _T_187; // @[Mux.scala 47:69]
  assign _GEN_15 = {{15'd0}, io_expected_out[9:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_189 = _GEN_15 << _T_188; // @[rawFloatFromFN.scala 54:36]
  assign _T_191 = {_T_189[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_16 = {{2'd0}, _T_188}; // @[rawFloatFromFN.scala 57:26]
  assign _T_192 = _GEN_16 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  assign _T_193 = _T_168 ? _T_192 : {{1'd0}, io_expected_out[14:10]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_194 = _T_168 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_17 = {{3'd0}, _T_194}; // @[rawFloatFromFN.scala 60:22]
  assign _T_195 = 5'h10 | _GEN_17; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_18 = {{1'd0}, _T_195}; // @[rawFloatFromFN.scala 59:15]
  assign _T_197 = _T_193 + _GEN_18; // @[rawFloatFromFN.scala 59:15]
  assign _T_198 = _T_168 & _T_169; // @[rawFloatFromFN.scala 62:34]
  assign _T_200 = _T_197[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_203 = _T_200 & ~_T_169; // @[rawFloatFromFN.scala 66:33]
  assign _T_206 = {1'b0,$signed(_T_197)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_208 = _T_168 ? _T_191 : io_expected_out[9:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_210 = {1'h0,~_T_198,_T_208}; // @[Cat.scala 29:58]
  assign _T_212 = _T_198 ? 3'h0 : _T_206[5:3]; // @[recFNFromFN.scala 48:16]
  assign _GEN_19 = {{2'd0}, _T_203}; // @[recFNFromFN.scala 48:79]
  assign _T_214 = _T_212 | _GEN_19; // @[recFNFromFN.scala 48:79]
  assign _T_217 = {_T_206[2:0],_T_210[9:0]}; // @[Cat.scala 29:58]
  assign _T_218 = {io_expected_out[15],_T_214}; // @[Cat.scala 29:58]
  assign _T_223 = io_actual_out[15:13] == 3'h0; // @[tests.scala 48:26]
  assign _T_225 = io_actual_out[15:13] == 3'h7; // @[tests.scala 48:55]
  assign _T_226 = _T_223 | _T_225; // @[tests.scala 48:39]
  assign _T_227 = io_actual_out[16:13] == io_expected_recOut[16:13]; // @[tests.scala 49:20]
  assign _T_230 = io_actual_out[9:0] == io_expected_recOut[9:0]; // @[tests.scala 49:54]
  assign _T_231 = _T_227 & _T_230; // @[tests.scala 49:31]
  assign _T_233 = io_actual_out[15:13] == 3'h6; // @[tests.scala 50:30]
  assign _T_235 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_236 = _T_233 ? _T_227 : _T_235; // @[tests.scala 50:16]
  assign _T_237 = _T_226 ? _T_231 : _T_236; // @[tests.scala 48:12]
  assign _T_238 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_MulAddRecFN.scala 82:35]
  assign io_expected_recOut = {_T_218,_T_217}; // @[ValExec_MulAddRecFN.scala 74:24]
  assign io_actual_out = mulAddRecFN_io_out; // @[ValExec_MulAddRecFN.scala 76:19]
  assign io_actual_exceptionFlags = mulAddRecFN_io_exceptionFlags; // @[ValExec_MulAddRecFN.scala 77:30]
  assign io_check = 1'h1; // @[ValExec_MulAddRecFN.scala 79:14]
  assign io_pass = _T_237 & _T_238; // @[ValExec_MulAddRecFN.scala 80:13]
  assign mulAddRecFN_io_a = {_T_53,_T_52}; // @[ValExec_MulAddRecFN.scala 68:22]
  assign mulAddRecFN_io_b = {_T_108,_T_107}; // @[ValExec_MulAddRecFN.scala 69:22]
  assign mulAddRecFN_io_c = {_T_163,_T_162}; // @[ValExec_MulAddRecFN.scala 70:22]
  assign mulAddRecFN_io_roundingMode = io_roundingMode; // @[ValExec_MulAddRecFN.scala 71:35]
  assign mulAddRecFN_io_detectTininess = io_detectTininess; // @[ValExec_MulAddRecFN.scala 72:35]
endmodule
