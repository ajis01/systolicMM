module CastFromNonLit(
  input  [6:0] io_in,
  output [6:0] io_out,
  output       io_valid
);
  wire  _T_2; // @[StrongEnum.scala 71:22]
  wire  _T_3; // @[StrongEnum.scala 71:22]
  wire  _T_4; // @[StrongEnum.scala 71:22]
  wire  _T_5; // @[StrongEnum.scala 71:22]
  wire  _T_6; // @[StrongEnum.scala 71:22]
  wire  _T_7; // @[StrongEnum.scala 71:22]
  wire  _T_8; // @[StrongEnum.scala 71:22]
  wire  _T_9; // @[StrongEnum.scala 71:22]
  assign _T_2 = io_out == 7'h0; // @[StrongEnum.scala 71:22]
  assign _T_3 = io_out == 7'h1; // @[StrongEnum.scala 71:22]
  assign _T_4 = io_out == 7'h2; // @[StrongEnum.scala 71:22]
  assign _T_5 = io_out == 7'h64; // @[StrongEnum.scala 71:22]
  assign _T_6 = io_out == 7'h65; // @[StrongEnum.scala 71:22]
  assign _T_7 = _T_2 | _T_3; // @[StrongEnum.scala 71:22]
  assign _T_8 = _T_7 | _T_4; // @[StrongEnum.scala 71:22]
  assign _T_9 = _T_8 | _T_5; // @[StrongEnum.scala 71:22]
  assign io_out = io_in; // @[StrongEnum.scala 70:10]
  assign io_valid = _T_9 | _T_6; // @[StrongEnum.scala 71:12]
endmodule
module CastFromNonLitTester(
  input   clock,
  input   reset
);
  wire [6:0] CastFromNonLit_io_in; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_io_out; // @[StrongEnum.scala 171:21]
  wire  CastFromNonLit_io_valid; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_1_io_in; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_1_io_out; // @[StrongEnum.scala 171:21]
  wire  CastFromNonLit_1_io_valid; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_2_io_in; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_2_io_out; // @[StrongEnum.scala 171:21]
  wire  CastFromNonLit_2_io_valid; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_3_io_in; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_3_io_out; // @[StrongEnum.scala 171:21]
  wire  CastFromNonLit_3_io_valid; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_4_io_in; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_4_io_out; // @[StrongEnum.scala 171:21]
  wire  CastFromNonLit_4_io_valid; // @[StrongEnum.scala 171:21]
  wire [6:0] CastFromNonLit_5_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_5_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_5_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_6_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_6_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_6_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_7_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_7_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_7_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_8_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_8_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_8_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_9_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_9_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_9_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_10_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_10_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_10_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_11_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_11_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_11_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_12_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_12_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_12_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_13_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_13_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_13_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_14_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_14_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_14_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_15_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_15_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_15_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_16_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_16_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_16_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_17_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_17_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_17_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_18_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_18_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_18_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_19_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_19_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_19_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_20_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_20_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_20_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_21_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_21_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_21_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_22_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_22_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_22_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_23_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_23_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_23_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_24_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_24_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_24_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_25_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_25_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_25_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_26_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_26_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_26_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_27_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_27_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_27_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_28_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_28_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_28_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_29_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_29_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_29_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_30_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_30_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_30_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_31_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_31_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_31_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_32_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_32_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_32_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_33_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_33_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_33_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_34_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_34_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_34_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_35_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_35_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_35_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_36_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_36_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_36_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_37_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_37_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_37_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_38_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_38_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_38_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_39_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_39_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_39_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_40_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_40_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_40_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_41_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_41_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_41_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_42_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_42_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_42_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_43_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_43_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_43_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_44_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_44_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_44_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_45_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_45_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_45_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_46_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_46_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_46_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_47_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_47_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_47_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_48_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_48_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_48_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_49_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_49_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_49_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_50_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_50_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_50_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_51_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_51_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_51_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_52_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_52_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_52_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_53_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_53_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_53_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_54_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_54_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_54_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_55_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_55_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_55_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_56_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_56_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_56_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_57_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_57_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_57_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_58_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_58_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_58_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_59_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_59_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_59_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_60_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_60_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_60_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_61_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_61_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_61_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_62_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_62_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_62_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_63_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_63_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_63_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_64_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_64_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_64_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_65_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_65_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_65_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_66_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_66_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_66_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_67_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_67_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_67_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_68_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_68_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_68_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_69_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_69_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_69_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_70_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_70_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_70_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_71_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_71_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_71_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_72_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_72_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_72_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_73_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_73_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_73_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_74_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_74_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_74_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_75_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_75_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_75_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_76_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_76_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_76_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_77_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_77_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_77_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_78_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_78_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_78_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_79_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_79_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_79_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_80_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_80_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_80_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_81_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_81_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_81_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_82_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_82_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_82_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_83_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_83_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_83_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_84_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_84_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_84_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_85_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_85_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_85_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_86_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_86_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_86_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_87_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_87_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_87_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_88_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_88_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_88_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_89_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_89_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_89_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_90_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_90_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_90_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_91_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_91_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_91_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_92_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_92_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_92_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_93_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_93_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_93_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_94_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_94_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_94_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_95_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_95_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_95_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_96_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_96_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_96_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_97_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_97_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_97_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_98_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_98_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_98_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_99_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_99_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_99_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_100_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_100_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_100_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_101_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_101_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_101_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_102_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_102_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_102_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_103_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_103_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_103_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_104_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_104_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_104_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_105_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_105_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_105_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_106_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_106_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_106_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_107_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_107_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_107_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_108_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_108_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_108_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_109_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_109_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_109_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_110_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_110_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_110_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_111_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_111_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_111_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_112_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_112_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_112_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_113_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_113_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_113_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_114_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_114_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_114_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_115_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_115_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_115_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_116_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_116_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_116_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_117_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_117_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_117_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_118_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_118_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_118_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_119_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_119_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_119_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_120_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_120_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_120_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_121_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_121_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_121_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_122_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_122_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_122_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_123_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_123_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_123_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_124_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_124_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_124_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_125_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_125_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_125_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_126_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_126_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_126_io_valid; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_127_io_in; // @[StrongEnum.scala 182:21]
  wire [6:0] CastFromNonLit_127_io_out; // @[StrongEnum.scala 182:21]
  wire  CastFromNonLit_127_io_valid; // @[StrongEnum.scala 182:21]
  wire  _T; // @[StrongEnum.scala 173:23]
  wire  _T_2; // @[StrongEnum.scala 173:11]
  wire  _T_3; // @[StrongEnum.scala 173:11]
  wire  _T_4; // @[StrongEnum.scala 174:25]
  wire  _T_6; // @[StrongEnum.scala 174:11]
  wire  _T_7; // @[StrongEnum.scala 174:11]
  wire  _T_8; // @[StrongEnum.scala 173:23]
  wire  _T_10; // @[StrongEnum.scala 173:11]
  wire  _T_11; // @[StrongEnum.scala 173:11]
  wire  _T_12; // @[StrongEnum.scala 174:25]
  wire  _T_14; // @[StrongEnum.scala 174:11]
  wire  _T_15; // @[StrongEnum.scala 174:11]
  wire  _T_16; // @[StrongEnum.scala 173:23]
  wire  _T_18; // @[StrongEnum.scala 173:11]
  wire  _T_19; // @[StrongEnum.scala 173:11]
  wire  _T_20; // @[StrongEnum.scala 174:25]
  wire  _T_22; // @[StrongEnum.scala 174:11]
  wire  _T_23; // @[StrongEnum.scala 174:11]
  wire  _T_24; // @[StrongEnum.scala 173:23]
  wire  _T_26; // @[StrongEnum.scala 173:11]
  wire  _T_27; // @[StrongEnum.scala 173:11]
  wire  _T_28; // @[StrongEnum.scala 174:25]
  wire  _T_30; // @[StrongEnum.scala 174:11]
  wire  _T_31; // @[StrongEnum.scala 174:11]
  wire  _T_32; // @[StrongEnum.scala 173:23]
  wire  _T_34; // @[StrongEnum.scala 173:11]
  wire  _T_35; // @[StrongEnum.scala 173:11]
  wire  _T_36; // @[StrongEnum.scala 174:25]
  wire  _T_38; // @[StrongEnum.scala 174:11]
  wire  _T_39; // @[StrongEnum.scala 174:11]
  wire  _T_40; // @[StrongEnum.scala 185:25]
  wire  _T_42; // @[StrongEnum.scala 185:11]
  wire  _T_43; // @[StrongEnum.scala 185:11]
  wire  _T_44; // @[StrongEnum.scala 185:25]
  wire  _T_46; // @[StrongEnum.scala 185:11]
  wire  _T_47; // @[StrongEnum.scala 185:11]
  wire  _T_48; // @[StrongEnum.scala 185:25]
  wire  _T_50; // @[StrongEnum.scala 185:11]
  wire  _T_51; // @[StrongEnum.scala 185:11]
  wire  _T_52; // @[StrongEnum.scala 185:25]
  wire  _T_54; // @[StrongEnum.scala 185:11]
  wire  _T_55; // @[StrongEnum.scala 185:11]
  wire  _T_56; // @[StrongEnum.scala 185:25]
  wire  _T_58; // @[StrongEnum.scala 185:11]
  wire  _T_59; // @[StrongEnum.scala 185:11]
  wire  _T_60; // @[StrongEnum.scala 185:25]
  wire  _T_62; // @[StrongEnum.scala 185:11]
  wire  _T_63; // @[StrongEnum.scala 185:11]
  wire  _T_64; // @[StrongEnum.scala 185:25]
  wire  _T_66; // @[StrongEnum.scala 185:11]
  wire  _T_67; // @[StrongEnum.scala 185:11]
  wire  _T_68; // @[StrongEnum.scala 185:25]
  wire  _T_70; // @[StrongEnum.scala 185:11]
  wire  _T_71; // @[StrongEnum.scala 185:11]
  wire  _T_72; // @[StrongEnum.scala 185:25]
  wire  _T_74; // @[StrongEnum.scala 185:11]
  wire  _T_75; // @[StrongEnum.scala 185:11]
  wire  _T_76; // @[StrongEnum.scala 185:25]
  wire  _T_78; // @[StrongEnum.scala 185:11]
  wire  _T_79; // @[StrongEnum.scala 185:11]
  wire  _T_80; // @[StrongEnum.scala 185:25]
  wire  _T_82; // @[StrongEnum.scala 185:11]
  wire  _T_83; // @[StrongEnum.scala 185:11]
  wire  _T_84; // @[StrongEnum.scala 185:25]
  wire  _T_86; // @[StrongEnum.scala 185:11]
  wire  _T_87; // @[StrongEnum.scala 185:11]
  wire  _T_88; // @[StrongEnum.scala 185:25]
  wire  _T_90; // @[StrongEnum.scala 185:11]
  wire  _T_91; // @[StrongEnum.scala 185:11]
  wire  _T_92; // @[StrongEnum.scala 185:25]
  wire  _T_94; // @[StrongEnum.scala 185:11]
  wire  _T_95; // @[StrongEnum.scala 185:11]
  wire  _T_96; // @[StrongEnum.scala 185:25]
  wire  _T_98; // @[StrongEnum.scala 185:11]
  wire  _T_99; // @[StrongEnum.scala 185:11]
  wire  _T_100; // @[StrongEnum.scala 185:25]
  wire  _T_102; // @[StrongEnum.scala 185:11]
  wire  _T_103; // @[StrongEnum.scala 185:11]
  wire  _T_104; // @[StrongEnum.scala 185:25]
  wire  _T_106; // @[StrongEnum.scala 185:11]
  wire  _T_107; // @[StrongEnum.scala 185:11]
  wire  _T_108; // @[StrongEnum.scala 185:25]
  wire  _T_110; // @[StrongEnum.scala 185:11]
  wire  _T_111; // @[StrongEnum.scala 185:11]
  wire  _T_112; // @[StrongEnum.scala 185:25]
  wire  _T_114; // @[StrongEnum.scala 185:11]
  wire  _T_115; // @[StrongEnum.scala 185:11]
  wire  _T_116; // @[StrongEnum.scala 185:25]
  wire  _T_118; // @[StrongEnum.scala 185:11]
  wire  _T_119; // @[StrongEnum.scala 185:11]
  wire  _T_120; // @[StrongEnum.scala 185:25]
  wire  _T_122; // @[StrongEnum.scala 185:11]
  wire  _T_123; // @[StrongEnum.scala 185:11]
  wire  _T_124; // @[StrongEnum.scala 185:25]
  wire  _T_126; // @[StrongEnum.scala 185:11]
  wire  _T_127; // @[StrongEnum.scala 185:11]
  wire  _T_128; // @[StrongEnum.scala 185:25]
  wire  _T_130; // @[StrongEnum.scala 185:11]
  wire  _T_131; // @[StrongEnum.scala 185:11]
  wire  _T_132; // @[StrongEnum.scala 185:25]
  wire  _T_134; // @[StrongEnum.scala 185:11]
  wire  _T_135; // @[StrongEnum.scala 185:11]
  wire  _T_136; // @[StrongEnum.scala 185:25]
  wire  _T_138; // @[StrongEnum.scala 185:11]
  wire  _T_139; // @[StrongEnum.scala 185:11]
  wire  _T_140; // @[StrongEnum.scala 185:25]
  wire  _T_142; // @[StrongEnum.scala 185:11]
  wire  _T_143; // @[StrongEnum.scala 185:11]
  wire  _T_144; // @[StrongEnum.scala 185:25]
  wire  _T_146; // @[StrongEnum.scala 185:11]
  wire  _T_147; // @[StrongEnum.scala 185:11]
  wire  _T_148; // @[StrongEnum.scala 185:25]
  wire  _T_150; // @[StrongEnum.scala 185:11]
  wire  _T_151; // @[StrongEnum.scala 185:11]
  wire  _T_152; // @[StrongEnum.scala 185:25]
  wire  _T_154; // @[StrongEnum.scala 185:11]
  wire  _T_155; // @[StrongEnum.scala 185:11]
  wire  _T_156; // @[StrongEnum.scala 185:25]
  wire  _T_158; // @[StrongEnum.scala 185:11]
  wire  _T_159; // @[StrongEnum.scala 185:11]
  wire  _T_160; // @[StrongEnum.scala 185:25]
  wire  _T_162; // @[StrongEnum.scala 185:11]
  wire  _T_163; // @[StrongEnum.scala 185:11]
  wire  _T_164; // @[StrongEnum.scala 185:25]
  wire  _T_166; // @[StrongEnum.scala 185:11]
  wire  _T_167; // @[StrongEnum.scala 185:11]
  wire  _T_168; // @[StrongEnum.scala 185:25]
  wire  _T_170; // @[StrongEnum.scala 185:11]
  wire  _T_171; // @[StrongEnum.scala 185:11]
  wire  _T_172; // @[StrongEnum.scala 185:25]
  wire  _T_174; // @[StrongEnum.scala 185:11]
  wire  _T_175; // @[StrongEnum.scala 185:11]
  wire  _T_176; // @[StrongEnum.scala 185:25]
  wire  _T_178; // @[StrongEnum.scala 185:11]
  wire  _T_179; // @[StrongEnum.scala 185:11]
  wire  _T_180; // @[StrongEnum.scala 185:25]
  wire  _T_182; // @[StrongEnum.scala 185:11]
  wire  _T_183; // @[StrongEnum.scala 185:11]
  wire  _T_184; // @[StrongEnum.scala 185:25]
  wire  _T_186; // @[StrongEnum.scala 185:11]
  wire  _T_187; // @[StrongEnum.scala 185:11]
  wire  _T_188; // @[StrongEnum.scala 185:25]
  wire  _T_190; // @[StrongEnum.scala 185:11]
  wire  _T_191; // @[StrongEnum.scala 185:11]
  wire  _T_192; // @[StrongEnum.scala 185:25]
  wire  _T_194; // @[StrongEnum.scala 185:11]
  wire  _T_195; // @[StrongEnum.scala 185:11]
  wire  _T_196; // @[StrongEnum.scala 185:25]
  wire  _T_198; // @[StrongEnum.scala 185:11]
  wire  _T_199; // @[StrongEnum.scala 185:11]
  wire  _T_200; // @[StrongEnum.scala 185:25]
  wire  _T_202; // @[StrongEnum.scala 185:11]
  wire  _T_203; // @[StrongEnum.scala 185:11]
  wire  _T_204; // @[StrongEnum.scala 185:25]
  wire  _T_206; // @[StrongEnum.scala 185:11]
  wire  _T_207; // @[StrongEnum.scala 185:11]
  wire  _T_208; // @[StrongEnum.scala 185:25]
  wire  _T_210; // @[StrongEnum.scala 185:11]
  wire  _T_211; // @[StrongEnum.scala 185:11]
  wire  _T_212; // @[StrongEnum.scala 185:25]
  wire  _T_214; // @[StrongEnum.scala 185:11]
  wire  _T_215; // @[StrongEnum.scala 185:11]
  wire  _T_216; // @[StrongEnum.scala 185:25]
  wire  _T_218; // @[StrongEnum.scala 185:11]
  wire  _T_219; // @[StrongEnum.scala 185:11]
  wire  _T_220; // @[StrongEnum.scala 185:25]
  wire  _T_222; // @[StrongEnum.scala 185:11]
  wire  _T_223; // @[StrongEnum.scala 185:11]
  wire  _T_224; // @[StrongEnum.scala 185:25]
  wire  _T_226; // @[StrongEnum.scala 185:11]
  wire  _T_227; // @[StrongEnum.scala 185:11]
  wire  _T_228; // @[StrongEnum.scala 185:25]
  wire  _T_230; // @[StrongEnum.scala 185:11]
  wire  _T_231; // @[StrongEnum.scala 185:11]
  wire  _T_232; // @[StrongEnum.scala 185:25]
  wire  _T_234; // @[StrongEnum.scala 185:11]
  wire  _T_235; // @[StrongEnum.scala 185:11]
  wire  _T_236; // @[StrongEnum.scala 185:25]
  wire  _T_238; // @[StrongEnum.scala 185:11]
  wire  _T_239; // @[StrongEnum.scala 185:11]
  wire  _T_240; // @[StrongEnum.scala 185:25]
  wire  _T_242; // @[StrongEnum.scala 185:11]
  wire  _T_243; // @[StrongEnum.scala 185:11]
  wire  _T_244; // @[StrongEnum.scala 185:25]
  wire  _T_246; // @[StrongEnum.scala 185:11]
  wire  _T_247; // @[StrongEnum.scala 185:11]
  wire  _T_248; // @[StrongEnum.scala 185:25]
  wire  _T_250; // @[StrongEnum.scala 185:11]
  wire  _T_251; // @[StrongEnum.scala 185:11]
  wire  _T_252; // @[StrongEnum.scala 185:25]
  wire  _T_254; // @[StrongEnum.scala 185:11]
  wire  _T_255; // @[StrongEnum.scala 185:11]
  wire  _T_256; // @[StrongEnum.scala 185:25]
  wire  _T_258; // @[StrongEnum.scala 185:11]
  wire  _T_259; // @[StrongEnum.scala 185:11]
  wire  _T_260; // @[StrongEnum.scala 185:25]
  wire  _T_262; // @[StrongEnum.scala 185:11]
  wire  _T_263; // @[StrongEnum.scala 185:11]
  wire  _T_264; // @[StrongEnum.scala 185:25]
  wire  _T_266; // @[StrongEnum.scala 185:11]
  wire  _T_267; // @[StrongEnum.scala 185:11]
  wire  _T_268; // @[StrongEnum.scala 185:25]
  wire  _T_270; // @[StrongEnum.scala 185:11]
  wire  _T_271; // @[StrongEnum.scala 185:11]
  wire  _T_272; // @[StrongEnum.scala 185:25]
  wire  _T_274; // @[StrongEnum.scala 185:11]
  wire  _T_275; // @[StrongEnum.scala 185:11]
  wire  _T_276; // @[StrongEnum.scala 185:25]
  wire  _T_278; // @[StrongEnum.scala 185:11]
  wire  _T_279; // @[StrongEnum.scala 185:11]
  wire  _T_280; // @[StrongEnum.scala 185:25]
  wire  _T_282; // @[StrongEnum.scala 185:11]
  wire  _T_283; // @[StrongEnum.scala 185:11]
  wire  _T_284; // @[StrongEnum.scala 185:25]
  wire  _T_286; // @[StrongEnum.scala 185:11]
  wire  _T_287; // @[StrongEnum.scala 185:11]
  wire  _T_288; // @[StrongEnum.scala 185:25]
  wire  _T_290; // @[StrongEnum.scala 185:11]
  wire  _T_291; // @[StrongEnum.scala 185:11]
  wire  _T_292; // @[StrongEnum.scala 185:25]
  wire  _T_294; // @[StrongEnum.scala 185:11]
  wire  _T_295; // @[StrongEnum.scala 185:11]
  wire  _T_296; // @[StrongEnum.scala 185:25]
  wire  _T_298; // @[StrongEnum.scala 185:11]
  wire  _T_299; // @[StrongEnum.scala 185:11]
  wire  _T_300; // @[StrongEnum.scala 185:25]
  wire  _T_302; // @[StrongEnum.scala 185:11]
  wire  _T_303; // @[StrongEnum.scala 185:11]
  wire  _T_304; // @[StrongEnum.scala 185:25]
  wire  _T_306; // @[StrongEnum.scala 185:11]
  wire  _T_307; // @[StrongEnum.scala 185:11]
  wire  _T_308; // @[StrongEnum.scala 185:25]
  wire  _T_310; // @[StrongEnum.scala 185:11]
  wire  _T_311; // @[StrongEnum.scala 185:11]
  wire  _T_312; // @[StrongEnum.scala 185:25]
  wire  _T_314; // @[StrongEnum.scala 185:11]
  wire  _T_315; // @[StrongEnum.scala 185:11]
  wire  _T_316; // @[StrongEnum.scala 185:25]
  wire  _T_318; // @[StrongEnum.scala 185:11]
  wire  _T_319; // @[StrongEnum.scala 185:11]
  wire  _T_320; // @[StrongEnum.scala 185:25]
  wire  _T_322; // @[StrongEnum.scala 185:11]
  wire  _T_323; // @[StrongEnum.scala 185:11]
  wire  _T_324; // @[StrongEnum.scala 185:25]
  wire  _T_326; // @[StrongEnum.scala 185:11]
  wire  _T_327; // @[StrongEnum.scala 185:11]
  wire  _T_328; // @[StrongEnum.scala 185:25]
  wire  _T_330; // @[StrongEnum.scala 185:11]
  wire  _T_331; // @[StrongEnum.scala 185:11]
  wire  _T_332; // @[StrongEnum.scala 185:25]
  wire  _T_334; // @[StrongEnum.scala 185:11]
  wire  _T_335; // @[StrongEnum.scala 185:11]
  wire  _T_336; // @[StrongEnum.scala 185:25]
  wire  _T_338; // @[StrongEnum.scala 185:11]
  wire  _T_339; // @[StrongEnum.scala 185:11]
  wire  _T_340; // @[StrongEnum.scala 185:25]
  wire  _T_342; // @[StrongEnum.scala 185:11]
  wire  _T_343; // @[StrongEnum.scala 185:11]
  wire  _T_344; // @[StrongEnum.scala 185:25]
  wire  _T_346; // @[StrongEnum.scala 185:11]
  wire  _T_347; // @[StrongEnum.scala 185:11]
  wire  _T_348; // @[StrongEnum.scala 185:25]
  wire  _T_350; // @[StrongEnum.scala 185:11]
  wire  _T_351; // @[StrongEnum.scala 185:11]
  wire  _T_352; // @[StrongEnum.scala 185:25]
  wire  _T_354; // @[StrongEnum.scala 185:11]
  wire  _T_355; // @[StrongEnum.scala 185:11]
  wire  _T_356; // @[StrongEnum.scala 185:25]
  wire  _T_358; // @[StrongEnum.scala 185:11]
  wire  _T_359; // @[StrongEnum.scala 185:11]
  wire  _T_360; // @[StrongEnum.scala 185:25]
  wire  _T_362; // @[StrongEnum.scala 185:11]
  wire  _T_363; // @[StrongEnum.scala 185:11]
  wire  _T_364; // @[StrongEnum.scala 185:25]
  wire  _T_366; // @[StrongEnum.scala 185:11]
  wire  _T_367; // @[StrongEnum.scala 185:11]
  wire  _T_368; // @[StrongEnum.scala 185:25]
  wire  _T_370; // @[StrongEnum.scala 185:11]
  wire  _T_371; // @[StrongEnum.scala 185:11]
  wire  _T_372; // @[StrongEnum.scala 185:25]
  wire  _T_374; // @[StrongEnum.scala 185:11]
  wire  _T_375; // @[StrongEnum.scala 185:11]
  wire  _T_376; // @[StrongEnum.scala 185:25]
  wire  _T_378; // @[StrongEnum.scala 185:11]
  wire  _T_379; // @[StrongEnum.scala 185:11]
  wire  _T_380; // @[StrongEnum.scala 185:25]
  wire  _T_382; // @[StrongEnum.scala 185:11]
  wire  _T_383; // @[StrongEnum.scala 185:11]
  wire  _T_384; // @[StrongEnum.scala 185:25]
  wire  _T_386; // @[StrongEnum.scala 185:11]
  wire  _T_387; // @[StrongEnum.scala 185:11]
  wire  _T_388; // @[StrongEnum.scala 185:25]
  wire  _T_390; // @[StrongEnum.scala 185:11]
  wire  _T_391; // @[StrongEnum.scala 185:11]
  wire  _T_392; // @[StrongEnum.scala 185:25]
  wire  _T_394; // @[StrongEnum.scala 185:11]
  wire  _T_395; // @[StrongEnum.scala 185:11]
  wire  _T_396; // @[StrongEnum.scala 185:25]
  wire  _T_398; // @[StrongEnum.scala 185:11]
  wire  _T_399; // @[StrongEnum.scala 185:11]
  wire  _T_400; // @[StrongEnum.scala 185:25]
  wire  _T_402; // @[StrongEnum.scala 185:11]
  wire  _T_403; // @[StrongEnum.scala 185:11]
  wire  _T_404; // @[StrongEnum.scala 185:25]
  wire  _T_406; // @[StrongEnum.scala 185:11]
  wire  _T_407; // @[StrongEnum.scala 185:11]
  wire  _T_408; // @[StrongEnum.scala 185:25]
  wire  _T_410; // @[StrongEnum.scala 185:11]
  wire  _T_411; // @[StrongEnum.scala 185:11]
  wire  _T_412; // @[StrongEnum.scala 185:25]
  wire  _T_414; // @[StrongEnum.scala 185:11]
  wire  _T_415; // @[StrongEnum.scala 185:11]
  wire  _T_416; // @[StrongEnum.scala 185:25]
  wire  _T_418; // @[StrongEnum.scala 185:11]
  wire  _T_419; // @[StrongEnum.scala 185:11]
  wire  _T_420; // @[StrongEnum.scala 185:25]
  wire  _T_422; // @[StrongEnum.scala 185:11]
  wire  _T_423; // @[StrongEnum.scala 185:11]
  wire  _T_424; // @[StrongEnum.scala 185:25]
  wire  _T_426; // @[StrongEnum.scala 185:11]
  wire  _T_427; // @[StrongEnum.scala 185:11]
  wire  _T_428; // @[StrongEnum.scala 185:25]
  wire  _T_430; // @[StrongEnum.scala 185:11]
  wire  _T_431; // @[StrongEnum.scala 185:11]
  wire  _T_432; // @[StrongEnum.scala 185:25]
  wire  _T_434; // @[StrongEnum.scala 185:11]
  wire  _T_435; // @[StrongEnum.scala 185:11]
  wire  _T_436; // @[StrongEnum.scala 185:25]
  wire  _T_438; // @[StrongEnum.scala 185:11]
  wire  _T_439; // @[StrongEnum.scala 185:11]
  wire  _T_440; // @[StrongEnum.scala 185:25]
  wire  _T_442; // @[StrongEnum.scala 185:11]
  wire  _T_443; // @[StrongEnum.scala 185:11]
  wire  _T_444; // @[StrongEnum.scala 185:25]
  wire  _T_446; // @[StrongEnum.scala 185:11]
  wire  _T_447; // @[StrongEnum.scala 185:11]
  wire  _T_448; // @[StrongEnum.scala 185:25]
  wire  _T_450; // @[StrongEnum.scala 185:11]
  wire  _T_451; // @[StrongEnum.scala 185:11]
  wire  _T_452; // @[StrongEnum.scala 185:25]
  wire  _T_454; // @[StrongEnum.scala 185:11]
  wire  _T_455; // @[StrongEnum.scala 185:11]
  wire  _T_456; // @[StrongEnum.scala 185:25]
  wire  _T_458; // @[StrongEnum.scala 185:11]
  wire  _T_459; // @[StrongEnum.scala 185:11]
  wire  _T_460; // @[StrongEnum.scala 185:25]
  wire  _T_462; // @[StrongEnum.scala 185:11]
  wire  _T_463; // @[StrongEnum.scala 185:11]
  wire  _T_464; // @[StrongEnum.scala 185:25]
  wire  _T_466; // @[StrongEnum.scala 185:11]
  wire  _T_467; // @[StrongEnum.scala 185:11]
  wire  _T_468; // @[StrongEnum.scala 185:25]
  wire  _T_470; // @[StrongEnum.scala 185:11]
  wire  _T_471; // @[StrongEnum.scala 185:11]
  wire  _T_472; // @[StrongEnum.scala 185:25]
  wire  _T_474; // @[StrongEnum.scala 185:11]
  wire  _T_475; // @[StrongEnum.scala 185:11]
  wire  _T_476; // @[StrongEnum.scala 185:25]
  wire  _T_478; // @[StrongEnum.scala 185:11]
  wire  _T_479; // @[StrongEnum.scala 185:11]
  wire  _T_480; // @[StrongEnum.scala 185:25]
  wire  _T_482; // @[StrongEnum.scala 185:11]
  wire  _T_483; // @[StrongEnum.scala 185:11]
  wire  _T_484; // @[StrongEnum.scala 185:25]
  wire  _T_486; // @[StrongEnum.scala 185:11]
  wire  _T_487; // @[StrongEnum.scala 185:11]
  wire  _T_488; // @[StrongEnum.scala 185:25]
  wire  _T_490; // @[StrongEnum.scala 185:11]
  wire  _T_491; // @[StrongEnum.scala 185:11]
  wire  _T_492; // @[StrongEnum.scala 185:25]
  wire  _T_494; // @[StrongEnum.scala 185:11]
  wire  _T_495; // @[StrongEnum.scala 185:11]
  wire  _T_496; // @[StrongEnum.scala 185:25]
  wire  _T_498; // @[StrongEnum.scala 185:11]
  wire  _T_499; // @[StrongEnum.scala 185:11]
  wire  _T_500; // @[StrongEnum.scala 185:25]
  wire  _T_502; // @[StrongEnum.scala 185:11]
  wire  _T_503; // @[StrongEnum.scala 185:11]
  wire  _T_504; // @[StrongEnum.scala 185:25]
  wire  _T_506; // @[StrongEnum.scala 185:11]
  wire  _T_507; // @[StrongEnum.scala 185:11]
  wire  _T_508; // @[StrongEnum.scala 185:25]
  wire  _T_510; // @[StrongEnum.scala 185:11]
  wire  _T_511; // @[StrongEnum.scala 185:11]
  wire  _T_512; // @[StrongEnum.scala 185:25]
  wire  _T_514; // @[StrongEnum.scala 185:11]
  wire  _T_515; // @[StrongEnum.scala 185:11]
  wire  _T_516; // @[StrongEnum.scala 185:25]
  wire  _T_518; // @[StrongEnum.scala 185:11]
  wire  _T_519; // @[StrongEnum.scala 185:11]
  wire  _T_520; // @[StrongEnum.scala 185:25]
  wire  _T_522; // @[StrongEnum.scala 185:11]
  wire  _T_523; // @[StrongEnum.scala 185:11]
  wire  _T_524; // @[StrongEnum.scala 185:25]
  wire  _T_526; // @[StrongEnum.scala 185:11]
  wire  _T_527; // @[StrongEnum.scala 185:11]
  wire  _T_528; // @[StrongEnum.scala 185:25]
  wire  _T_530; // @[StrongEnum.scala 185:11]
  wire  _T_531; // @[StrongEnum.scala 185:11]
  wire  _T_533; // @[StrongEnum.scala 188:7]
  CastFromNonLit CastFromNonLit ( // @[StrongEnum.scala 171:21]
    .io_in(CastFromNonLit_io_in),
    .io_out(CastFromNonLit_io_out),
    .io_valid(CastFromNonLit_io_valid)
  );
  CastFromNonLit CastFromNonLit_1 ( // @[StrongEnum.scala 171:21]
    .io_in(CastFromNonLit_1_io_in),
    .io_out(CastFromNonLit_1_io_out),
    .io_valid(CastFromNonLit_1_io_valid)
  );
  CastFromNonLit CastFromNonLit_2 ( // @[StrongEnum.scala 171:21]
    .io_in(CastFromNonLit_2_io_in),
    .io_out(CastFromNonLit_2_io_out),
    .io_valid(CastFromNonLit_2_io_valid)
  );
  CastFromNonLit CastFromNonLit_3 ( // @[StrongEnum.scala 171:21]
    .io_in(CastFromNonLit_3_io_in),
    .io_out(CastFromNonLit_3_io_out),
    .io_valid(CastFromNonLit_3_io_valid)
  );
  CastFromNonLit CastFromNonLit_4 ( // @[StrongEnum.scala 171:21]
    .io_in(CastFromNonLit_4_io_in),
    .io_out(CastFromNonLit_4_io_out),
    .io_valid(CastFromNonLit_4_io_valid)
  );
  CastFromNonLit CastFromNonLit_5 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_5_io_in),
    .io_out(CastFromNonLit_5_io_out),
    .io_valid(CastFromNonLit_5_io_valid)
  );
  CastFromNonLit CastFromNonLit_6 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_6_io_in),
    .io_out(CastFromNonLit_6_io_out),
    .io_valid(CastFromNonLit_6_io_valid)
  );
  CastFromNonLit CastFromNonLit_7 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_7_io_in),
    .io_out(CastFromNonLit_7_io_out),
    .io_valid(CastFromNonLit_7_io_valid)
  );
  CastFromNonLit CastFromNonLit_8 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_8_io_in),
    .io_out(CastFromNonLit_8_io_out),
    .io_valid(CastFromNonLit_8_io_valid)
  );
  CastFromNonLit CastFromNonLit_9 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_9_io_in),
    .io_out(CastFromNonLit_9_io_out),
    .io_valid(CastFromNonLit_9_io_valid)
  );
  CastFromNonLit CastFromNonLit_10 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_10_io_in),
    .io_out(CastFromNonLit_10_io_out),
    .io_valid(CastFromNonLit_10_io_valid)
  );
  CastFromNonLit CastFromNonLit_11 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_11_io_in),
    .io_out(CastFromNonLit_11_io_out),
    .io_valid(CastFromNonLit_11_io_valid)
  );
  CastFromNonLit CastFromNonLit_12 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_12_io_in),
    .io_out(CastFromNonLit_12_io_out),
    .io_valid(CastFromNonLit_12_io_valid)
  );
  CastFromNonLit CastFromNonLit_13 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_13_io_in),
    .io_out(CastFromNonLit_13_io_out),
    .io_valid(CastFromNonLit_13_io_valid)
  );
  CastFromNonLit CastFromNonLit_14 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_14_io_in),
    .io_out(CastFromNonLit_14_io_out),
    .io_valid(CastFromNonLit_14_io_valid)
  );
  CastFromNonLit CastFromNonLit_15 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_15_io_in),
    .io_out(CastFromNonLit_15_io_out),
    .io_valid(CastFromNonLit_15_io_valid)
  );
  CastFromNonLit CastFromNonLit_16 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_16_io_in),
    .io_out(CastFromNonLit_16_io_out),
    .io_valid(CastFromNonLit_16_io_valid)
  );
  CastFromNonLit CastFromNonLit_17 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_17_io_in),
    .io_out(CastFromNonLit_17_io_out),
    .io_valid(CastFromNonLit_17_io_valid)
  );
  CastFromNonLit CastFromNonLit_18 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_18_io_in),
    .io_out(CastFromNonLit_18_io_out),
    .io_valid(CastFromNonLit_18_io_valid)
  );
  CastFromNonLit CastFromNonLit_19 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_19_io_in),
    .io_out(CastFromNonLit_19_io_out),
    .io_valid(CastFromNonLit_19_io_valid)
  );
  CastFromNonLit CastFromNonLit_20 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_20_io_in),
    .io_out(CastFromNonLit_20_io_out),
    .io_valid(CastFromNonLit_20_io_valid)
  );
  CastFromNonLit CastFromNonLit_21 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_21_io_in),
    .io_out(CastFromNonLit_21_io_out),
    .io_valid(CastFromNonLit_21_io_valid)
  );
  CastFromNonLit CastFromNonLit_22 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_22_io_in),
    .io_out(CastFromNonLit_22_io_out),
    .io_valid(CastFromNonLit_22_io_valid)
  );
  CastFromNonLit CastFromNonLit_23 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_23_io_in),
    .io_out(CastFromNonLit_23_io_out),
    .io_valid(CastFromNonLit_23_io_valid)
  );
  CastFromNonLit CastFromNonLit_24 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_24_io_in),
    .io_out(CastFromNonLit_24_io_out),
    .io_valid(CastFromNonLit_24_io_valid)
  );
  CastFromNonLit CastFromNonLit_25 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_25_io_in),
    .io_out(CastFromNonLit_25_io_out),
    .io_valid(CastFromNonLit_25_io_valid)
  );
  CastFromNonLit CastFromNonLit_26 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_26_io_in),
    .io_out(CastFromNonLit_26_io_out),
    .io_valid(CastFromNonLit_26_io_valid)
  );
  CastFromNonLit CastFromNonLit_27 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_27_io_in),
    .io_out(CastFromNonLit_27_io_out),
    .io_valid(CastFromNonLit_27_io_valid)
  );
  CastFromNonLit CastFromNonLit_28 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_28_io_in),
    .io_out(CastFromNonLit_28_io_out),
    .io_valid(CastFromNonLit_28_io_valid)
  );
  CastFromNonLit CastFromNonLit_29 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_29_io_in),
    .io_out(CastFromNonLit_29_io_out),
    .io_valid(CastFromNonLit_29_io_valid)
  );
  CastFromNonLit CastFromNonLit_30 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_30_io_in),
    .io_out(CastFromNonLit_30_io_out),
    .io_valid(CastFromNonLit_30_io_valid)
  );
  CastFromNonLit CastFromNonLit_31 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_31_io_in),
    .io_out(CastFromNonLit_31_io_out),
    .io_valid(CastFromNonLit_31_io_valid)
  );
  CastFromNonLit CastFromNonLit_32 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_32_io_in),
    .io_out(CastFromNonLit_32_io_out),
    .io_valid(CastFromNonLit_32_io_valid)
  );
  CastFromNonLit CastFromNonLit_33 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_33_io_in),
    .io_out(CastFromNonLit_33_io_out),
    .io_valid(CastFromNonLit_33_io_valid)
  );
  CastFromNonLit CastFromNonLit_34 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_34_io_in),
    .io_out(CastFromNonLit_34_io_out),
    .io_valid(CastFromNonLit_34_io_valid)
  );
  CastFromNonLit CastFromNonLit_35 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_35_io_in),
    .io_out(CastFromNonLit_35_io_out),
    .io_valid(CastFromNonLit_35_io_valid)
  );
  CastFromNonLit CastFromNonLit_36 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_36_io_in),
    .io_out(CastFromNonLit_36_io_out),
    .io_valid(CastFromNonLit_36_io_valid)
  );
  CastFromNonLit CastFromNonLit_37 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_37_io_in),
    .io_out(CastFromNonLit_37_io_out),
    .io_valid(CastFromNonLit_37_io_valid)
  );
  CastFromNonLit CastFromNonLit_38 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_38_io_in),
    .io_out(CastFromNonLit_38_io_out),
    .io_valid(CastFromNonLit_38_io_valid)
  );
  CastFromNonLit CastFromNonLit_39 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_39_io_in),
    .io_out(CastFromNonLit_39_io_out),
    .io_valid(CastFromNonLit_39_io_valid)
  );
  CastFromNonLit CastFromNonLit_40 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_40_io_in),
    .io_out(CastFromNonLit_40_io_out),
    .io_valid(CastFromNonLit_40_io_valid)
  );
  CastFromNonLit CastFromNonLit_41 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_41_io_in),
    .io_out(CastFromNonLit_41_io_out),
    .io_valid(CastFromNonLit_41_io_valid)
  );
  CastFromNonLit CastFromNonLit_42 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_42_io_in),
    .io_out(CastFromNonLit_42_io_out),
    .io_valid(CastFromNonLit_42_io_valid)
  );
  CastFromNonLit CastFromNonLit_43 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_43_io_in),
    .io_out(CastFromNonLit_43_io_out),
    .io_valid(CastFromNonLit_43_io_valid)
  );
  CastFromNonLit CastFromNonLit_44 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_44_io_in),
    .io_out(CastFromNonLit_44_io_out),
    .io_valid(CastFromNonLit_44_io_valid)
  );
  CastFromNonLit CastFromNonLit_45 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_45_io_in),
    .io_out(CastFromNonLit_45_io_out),
    .io_valid(CastFromNonLit_45_io_valid)
  );
  CastFromNonLit CastFromNonLit_46 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_46_io_in),
    .io_out(CastFromNonLit_46_io_out),
    .io_valid(CastFromNonLit_46_io_valid)
  );
  CastFromNonLit CastFromNonLit_47 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_47_io_in),
    .io_out(CastFromNonLit_47_io_out),
    .io_valid(CastFromNonLit_47_io_valid)
  );
  CastFromNonLit CastFromNonLit_48 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_48_io_in),
    .io_out(CastFromNonLit_48_io_out),
    .io_valid(CastFromNonLit_48_io_valid)
  );
  CastFromNonLit CastFromNonLit_49 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_49_io_in),
    .io_out(CastFromNonLit_49_io_out),
    .io_valid(CastFromNonLit_49_io_valid)
  );
  CastFromNonLit CastFromNonLit_50 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_50_io_in),
    .io_out(CastFromNonLit_50_io_out),
    .io_valid(CastFromNonLit_50_io_valid)
  );
  CastFromNonLit CastFromNonLit_51 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_51_io_in),
    .io_out(CastFromNonLit_51_io_out),
    .io_valid(CastFromNonLit_51_io_valid)
  );
  CastFromNonLit CastFromNonLit_52 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_52_io_in),
    .io_out(CastFromNonLit_52_io_out),
    .io_valid(CastFromNonLit_52_io_valid)
  );
  CastFromNonLit CastFromNonLit_53 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_53_io_in),
    .io_out(CastFromNonLit_53_io_out),
    .io_valid(CastFromNonLit_53_io_valid)
  );
  CastFromNonLit CastFromNonLit_54 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_54_io_in),
    .io_out(CastFromNonLit_54_io_out),
    .io_valid(CastFromNonLit_54_io_valid)
  );
  CastFromNonLit CastFromNonLit_55 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_55_io_in),
    .io_out(CastFromNonLit_55_io_out),
    .io_valid(CastFromNonLit_55_io_valid)
  );
  CastFromNonLit CastFromNonLit_56 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_56_io_in),
    .io_out(CastFromNonLit_56_io_out),
    .io_valid(CastFromNonLit_56_io_valid)
  );
  CastFromNonLit CastFromNonLit_57 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_57_io_in),
    .io_out(CastFromNonLit_57_io_out),
    .io_valid(CastFromNonLit_57_io_valid)
  );
  CastFromNonLit CastFromNonLit_58 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_58_io_in),
    .io_out(CastFromNonLit_58_io_out),
    .io_valid(CastFromNonLit_58_io_valid)
  );
  CastFromNonLit CastFromNonLit_59 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_59_io_in),
    .io_out(CastFromNonLit_59_io_out),
    .io_valid(CastFromNonLit_59_io_valid)
  );
  CastFromNonLit CastFromNonLit_60 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_60_io_in),
    .io_out(CastFromNonLit_60_io_out),
    .io_valid(CastFromNonLit_60_io_valid)
  );
  CastFromNonLit CastFromNonLit_61 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_61_io_in),
    .io_out(CastFromNonLit_61_io_out),
    .io_valid(CastFromNonLit_61_io_valid)
  );
  CastFromNonLit CastFromNonLit_62 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_62_io_in),
    .io_out(CastFromNonLit_62_io_out),
    .io_valid(CastFromNonLit_62_io_valid)
  );
  CastFromNonLit CastFromNonLit_63 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_63_io_in),
    .io_out(CastFromNonLit_63_io_out),
    .io_valid(CastFromNonLit_63_io_valid)
  );
  CastFromNonLit CastFromNonLit_64 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_64_io_in),
    .io_out(CastFromNonLit_64_io_out),
    .io_valid(CastFromNonLit_64_io_valid)
  );
  CastFromNonLit CastFromNonLit_65 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_65_io_in),
    .io_out(CastFromNonLit_65_io_out),
    .io_valid(CastFromNonLit_65_io_valid)
  );
  CastFromNonLit CastFromNonLit_66 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_66_io_in),
    .io_out(CastFromNonLit_66_io_out),
    .io_valid(CastFromNonLit_66_io_valid)
  );
  CastFromNonLit CastFromNonLit_67 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_67_io_in),
    .io_out(CastFromNonLit_67_io_out),
    .io_valid(CastFromNonLit_67_io_valid)
  );
  CastFromNonLit CastFromNonLit_68 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_68_io_in),
    .io_out(CastFromNonLit_68_io_out),
    .io_valid(CastFromNonLit_68_io_valid)
  );
  CastFromNonLit CastFromNonLit_69 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_69_io_in),
    .io_out(CastFromNonLit_69_io_out),
    .io_valid(CastFromNonLit_69_io_valid)
  );
  CastFromNonLit CastFromNonLit_70 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_70_io_in),
    .io_out(CastFromNonLit_70_io_out),
    .io_valid(CastFromNonLit_70_io_valid)
  );
  CastFromNonLit CastFromNonLit_71 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_71_io_in),
    .io_out(CastFromNonLit_71_io_out),
    .io_valid(CastFromNonLit_71_io_valid)
  );
  CastFromNonLit CastFromNonLit_72 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_72_io_in),
    .io_out(CastFromNonLit_72_io_out),
    .io_valid(CastFromNonLit_72_io_valid)
  );
  CastFromNonLit CastFromNonLit_73 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_73_io_in),
    .io_out(CastFromNonLit_73_io_out),
    .io_valid(CastFromNonLit_73_io_valid)
  );
  CastFromNonLit CastFromNonLit_74 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_74_io_in),
    .io_out(CastFromNonLit_74_io_out),
    .io_valid(CastFromNonLit_74_io_valid)
  );
  CastFromNonLit CastFromNonLit_75 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_75_io_in),
    .io_out(CastFromNonLit_75_io_out),
    .io_valid(CastFromNonLit_75_io_valid)
  );
  CastFromNonLit CastFromNonLit_76 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_76_io_in),
    .io_out(CastFromNonLit_76_io_out),
    .io_valid(CastFromNonLit_76_io_valid)
  );
  CastFromNonLit CastFromNonLit_77 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_77_io_in),
    .io_out(CastFromNonLit_77_io_out),
    .io_valid(CastFromNonLit_77_io_valid)
  );
  CastFromNonLit CastFromNonLit_78 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_78_io_in),
    .io_out(CastFromNonLit_78_io_out),
    .io_valid(CastFromNonLit_78_io_valid)
  );
  CastFromNonLit CastFromNonLit_79 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_79_io_in),
    .io_out(CastFromNonLit_79_io_out),
    .io_valid(CastFromNonLit_79_io_valid)
  );
  CastFromNonLit CastFromNonLit_80 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_80_io_in),
    .io_out(CastFromNonLit_80_io_out),
    .io_valid(CastFromNonLit_80_io_valid)
  );
  CastFromNonLit CastFromNonLit_81 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_81_io_in),
    .io_out(CastFromNonLit_81_io_out),
    .io_valid(CastFromNonLit_81_io_valid)
  );
  CastFromNonLit CastFromNonLit_82 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_82_io_in),
    .io_out(CastFromNonLit_82_io_out),
    .io_valid(CastFromNonLit_82_io_valid)
  );
  CastFromNonLit CastFromNonLit_83 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_83_io_in),
    .io_out(CastFromNonLit_83_io_out),
    .io_valid(CastFromNonLit_83_io_valid)
  );
  CastFromNonLit CastFromNonLit_84 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_84_io_in),
    .io_out(CastFromNonLit_84_io_out),
    .io_valid(CastFromNonLit_84_io_valid)
  );
  CastFromNonLit CastFromNonLit_85 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_85_io_in),
    .io_out(CastFromNonLit_85_io_out),
    .io_valid(CastFromNonLit_85_io_valid)
  );
  CastFromNonLit CastFromNonLit_86 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_86_io_in),
    .io_out(CastFromNonLit_86_io_out),
    .io_valid(CastFromNonLit_86_io_valid)
  );
  CastFromNonLit CastFromNonLit_87 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_87_io_in),
    .io_out(CastFromNonLit_87_io_out),
    .io_valid(CastFromNonLit_87_io_valid)
  );
  CastFromNonLit CastFromNonLit_88 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_88_io_in),
    .io_out(CastFromNonLit_88_io_out),
    .io_valid(CastFromNonLit_88_io_valid)
  );
  CastFromNonLit CastFromNonLit_89 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_89_io_in),
    .io_out(CastFromNonLit_89_io_out),
    .io_valid(CastFromNonLit_89_io_valid)
  );
  CastFromNonLit CastFromNonLit_90 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_90_io_in),
    .io_out(CastFromNonLit_90_io_out),
    .io_valid(CastFromNonLit_90_io_valid)
  );
  CastFromNonLit CastFromNonLit_91 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_91_io_in),
    .io_out(CastFromNonLit_91_io_out),
    .io_valid(CastFromNonLit_91_io_valid)
  );
  CastFromNonLit CastFromNonLit_92 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_92_io_in),
    .io_out(CastFromNonLit_92_io_out),
    .io_valid(CastFromNonLit_92_io_valid)
  );
  CastFromNonLit CastFromNonLit_93 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_93_io_in),
    .io_out(CastFromNonLit_93_io_out),
    .io_valid(CastFromNonLit_93_io_valid)
  );
  CastFromNonLit CastFromNonLit_94 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_94_io_in),
    .io_out(CastFromNonLit_94_io_out),
    .io_valid(CastFromNonLit_94_io_valid)
  );
  CastFromNonLit CastFromNonLit_95 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_95_io_in),
    .io_out(CastFromNonLit_95_io_out),
    .io_valid(CastFromNonLit_95_io_valid)
  );
  CastFromNonLit CastFromNonLit_96 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_96_io_in),
    .io_out(CastFromNonLit_96_io_out),
    .io_valid(CastFromNonLit_96_io_valid)
  );
  CastFromNonLit CastFromNonLit_97 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_97_io_in),
    .io_out(CastFromNonLit_97_io_out),
    .io_valid(CastFromNonLit_97_io_valid)
  );
  CastFromNonLit CastFromNonLit_98 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_98_io_in),
    .io_out(CastFromNonLit_98_io_out),
    .io_valid(CastFromNonLit_98_io_valid)
  );
  CastFromNonLit CastFromNonLit_99 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_99_io_in),
    .io_out(CastFromNonLit_99_io_out),
    .io_valid(CastFromNonLit_99_io_valid)
  );
  CastFromNonLit CastFromNonLit_100 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_100_io_in),
    .io_out(CastFromNonLit_100_io_out),
    .io_valid(CastFromNonLit_100_io_valid)
  );
  CastFromNonLit CastFromNonLit_101 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_101_io_in),
    .io_out(CastFromNonLit_101_io_out),
    .io_valid(CastFromNonLit_101_io_valid)
  );
  CastFromNonLit CastFromNonLit_102 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_102_io_in),
    .io_out(CastFromNonLit_102_io_out),
    .io_valid(CastFromNonLit_102_io_valid)
  );
  CastFromNonLit CastFromNonLit_103 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_103_io_in),
    .io_out(CastFromNonLit_103_io_out),
    .io_valid(CastFromNonLit_103_io_valid)
  );
  CastFromNonLit CastFromNonLit_104 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_104_io_in),
    .io_out(CastFromNonLit_104_io_out),
    .io_valid(CastFromNonLit_104_io_valid)
  );
  CastFromNonLit CastFromNonLit_105 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_105_io_in),
    .io_out(CastFromNonLit_105_io_out),
    .io_valid(CastFromNonLit_105_io_valid)
  );
  CastFromNonLit CastFromNonLit_106 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_106_io_in),
    .io_out(CastFromNonLit_106_io_out),
    .io_valid(CastFromNonLit_106_io_valid)
  );
  CastFromNonLit CastFromNonLit_107 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_107_io_in),
    .io_out(CastFromNonLit_107_io_out),
    .io_valid(CastFromNonLit_107_io_valid)
  );
  CastFromNonLit CastFromNonLit_108 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_108_io_in),
    .io_out(CastFromNonLit_108_io_out),
    .io_valid(CastFromNonLit_108_io_valid)
  );
  CastFromNonLit CastFromNonLit_109 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_109_io_in),
    .io_out(CastFromNonLit_109_io_out),
    .io_valid(CastFromNonLit_109_io_valid)
  );
  CastFromNonLit CastFromNonLit_110 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_110_io_in),
    .io_out(CastFromNonLit_110_io_out),
    .io_valid(CastFromNonLit_110_io_valid)
  );
  CastFromNonLit CastFromNonLit_111 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_111_io_in),
    .io_out(CastFromNonLit_111_io_out),
    .io_valid(CastFromNonLit_111_io_valid)
  );
  CastFromNonLit CastFromNonLit_112 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_112_io_in),
    .io_out(CastFromNonLit_112_io_out),
    .io_valid(CastFromNonLit_112_io_valid)
  );
  CastFromNonLit CastFromNonLit_113 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_113_io_in),
    .io_out(CastFromNonLit_113_io_out),
    .io_valid(CastFromNonLit_113_io_valid)
  );
  CastFromNonLit CastFromNonLit_114 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_114_io_in),
    .io_out(CastFromNonLit_114_io_out),
    .io_valid(CastFromNonLit_114_io_valid)
  );
  CastFromNonLit CastFromNonLit_115 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_115_io_in),
    .io_out(CastFromNonLit_115_io_out),
    .io_valid(CastFromNonLit_115_io_valid)
  );
  CastFromNonLit CastFromNonLit_116 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_116_io_in),
    .io_out(CastFromNonLit_116_io_out),
    .io_valid(CastFromNonLit_116_io_valid)
  );
  CastFromNonLit CastFromNonLit_117 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_117_io_in),
    .io_out(CastFromNonLit_117_io_out),
    .io_valid(CastFromNonLit_117_io_valid)
  );
  CastFromNonLit CastFromNonLit_118 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_118_io_in),
    .io_out(CastFromNonLit_118_io_out),
    .io_valid(CastFromNonLit_118_io_valid)
  );
  CastFromNonLit CastFromNonLit_119 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_119_io_in),
    .io_out(CastFromNonLit_119_io_out),
    .io_valid(CastFromNonLit_119_io_valid)
  );
  CastFromNonLit CastFromNonLit_120 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_120_io_in),
    .io_out(CastFromNonLit_120_io_out),
    .io_valid(CastFromNonLit_120_io_valid)
  );
  CastFromNonLit CastFromNonLit_121 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_121_io_in),
    .io_out(CastFromNonLit_121_io_out),
    .io_valid(CastFromNonLit_121_io_valid)
  );
  CastFromNonLit CastFromNonLit_122 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_122_io_in),
    .io_out(CastFromNonLit_122_io_out),
    .io_valid(CastFromNonLit_122_io_valid)
  );
  CastFromNonLit CastFromNonLit_123 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_123_io_in),
    .io_out(CastFromNonLit_123_io_out),
    .io_valid(CastFromNonLit_123_io_valid)
  );
  CastFromNonLit CastFromNonLit_124 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_124_io_in),
    .io_out(CastFromNonLit_124_io_out),
    .io_valid(CastFromNonLit_124_io_valid)
  );
  CastFromNonLit CastFromNonLit_125 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_125_io_in),
    .io_out(CastFromNonLit_125_io_out),
    .io_valid(CastFromNonLit_125_io_valid)
  );
  CastFromNonLit CastFromNonLit_126 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_126_io_in),
    .io_out(CastFromNonLit_126_io_out),
    .io_valid(CastFromNonLit_126_io_valid)
  );
  CastFromNonLit CastFromNonLit_127 ( // @[StrongEnum.scala 182:21]
    .io_in(CastFromNonLit_127_io_in),
    .io_out(CastFromNonLit_127_io_out),
    .io_valid(CastFromNonLit_127_io_valid)
  );
  assign _T = CastFromNonLit_io_out == 7'h0; // @[StrongEnum.scala 173:23]
  assign _T_2 = _T | reset; // @[StrongEnum.scala 173:11]
  assign _T_3 = _T_2 == 1'h0; // @[StrongEnum.scala 173:11]
  assign _T_4 = CastFromNonLit_io_valid; // @[StrongEnum.scala 174:25]
  assign _T_6 = _T_4 | reset; // @[StrongEnum.scala 174:11]
  assign _T_7 = _T_6 == 1'h0; // @[StrongEnum.scala 174:11]
  assign _T_8 = CastFromNonLit_1_io_out == 7'h1; // @[StrongEnum.scala 173:23]
  assign _T_10 = _T_8 | reset; // @[StrongEnum.scala 173:11]
  assign _T_11 = _T_10 == 1'h0; // @[StrongEnum.scala 173:11]
  assign _T_12 = CastFromNonLit_1_io_valid; // @[StrongEnum.scala 174:25]
  assign _T_14 = _T_12 | reset; // @[StrongEnum.scala 174:11]
  assign _T_15 = _T_14 == 1'h0; // @[StrongEnum.scala 174:11]
  assign _T_16 = CastFromNonLit_2_io_out == 7'h2; // @[StrongEnum.scala 173:23]
  assign _T_18 = _T_16 | reset; // @[StrongEnum.scala 173:11]
  assign _T_19 = _T_18 == 1'h0; // @[StrongEnum.scala 173:11]
  assign _T_20 = CastFromNonLit_2_io_valid; // @[StrongEnum.scala 174:25]
  assign _T_22 = _T_20 | reset; // @[StrongEnum.scala 174:11]
  assign _T_23 = _T_22 == 1'h0; // @[StrongEnum.scala 174:11]
  assign _T_24 = CastFromNonLit_3_io_out == 7'h64; // @[StrongEnum.scala 173:23]
  assign _T_26 = _T_24 | reset; // @[StrongEnum.scala 173:11]
  assign _T_27 = _T_26 == 1'h0; // @[StrongEnum.scala 173:11]
  assign _T_28 = CastFromNonLit_3_io_valid; // @[StrongEnum.scala 174:25]
  assign _T_30 = _T_28 | reset; // @[StrongEnum.scala 174:11]
  assign _T_31 = _T_30 == 1'h0; // @[StrongEnum.scala 174:11]
  assign _T_32 = CastFromNonLit_4_io_out == 7'h65; // @[StrongEnum.scala 173:23]
  assign _T_34 = _T_32 | reset; // @[StrongEnum.scala 173:11]
  assign _T_35 = _T_34 == 1'h0; // @[StrongEnum.scala 173:11]
  assign _T_36 = CastFromNonLit_4_io_valid; // @[StrongEnum.scala 174:25]
  assign _T_38 = _T_36 | reset; // @[StrongEnum.scala 174:11]
  assign _T_39 = _T_38 == 1'h0; // @[StrongEnum.scala 174:11]
  assign _T_40 = CastFromNonLit_5_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_42 = _T_40 | reset; // @[StrongEnum.scala 185:11]
  assign _T_43 = _T_42 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_44 = CastFromNonLit_6_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_46 = _T_44 | reset; // @[StrongEnum.scala 185:11]
  assign _T_47 = _T_46 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_48 = CastFromNonLit_7_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_50 = _T_48 | reset; // @[StrongEnum.scala 185:11]
  assign _T_51 = _T_50 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_52 = CastFromNonLit_8_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_54 = _T_52 | reset; // @[StrongEnum.scala 185:11]
  assign _T_55 = _T_54 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_56 = CastFromNonLit_9_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_58 = _T_56 | reset; // @[StrongEnum.scala 185:11]
  assign _T_59 = _T_58 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_60 = CastFromNonLit_10_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_62 = _T_60 | reset; // @[StrongEnum.scala 185:11]
  assign _T_63 = _T_62 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_64 = CastFromNonLit_11_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_66 = _T_64 | reset; // @[StrongEnum.scala 185:11]
  assign _T_67 = _T_66 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_68 = CastFromNonLit_12_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_70 = _T_68 | reset; // @[StrongEnum.scala 185:11]
  assign _T_71 = _T_70 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_72 = CastFromNonLit_13_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_74 = _T_72 | reset; // @[StrongEnum.scala 185:11]
  assign _T_75 = _T_74 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_76 = CastFromNonLit_14_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_78 = _T_76 | reset; // @[StrongEnum.scala 185:11]
  assign _T_79 = _T_78 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_80 = CastFromNonLit_15_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_82 = _T_80 | reset; // @[StrongEnum.scala 185:11]
  assign _T_83 = _T_82 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_84 = CastFromNonLit_16_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_86 = _T_84 | reset; // @[StrongEnum.scala 185:11]
  assign _T_87 = _T_86 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_88 = CastFromNonLit_17_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_90 = _T_88 | reset; // @[StrongEnum.scala 185:11]
  assign _T_91 = _T_90 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_92 = CastFromNonLit_18_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_94 = _T_92 | reset; // @[StrongEnum.scala 185:11]
  assign _T_95 = _T_94 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_96 = CastFromNonLit_19_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_98 = _T_96 | reset; // @[StrongEnum.scala 185:11]
  assign _T_99 = _T_98 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_100 = CastFromNonLit_20_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_102 = _T_100 | reset; // @[StrongEnum.scala 185:11]
  assign _T_103 = _T_102 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_104 = CastFromNonLit_21_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_106 = _T_104 | reset; // @[StrongEnum.scala 185:11]
  assign _T_107 = _T_106 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_108 = CastFromNonLit_22_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_110 = _T_108 | reset; // @[StrongEnum.scala 185:11]
  assign _T_111 = _T_110 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_112 = CastFromNonLit_23_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_114 = _T_112 | reset; // @[StrongEnum.scala 185:11]
  assign _T_115 = _T_114 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_116 = CastFromNonLit_24_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_118 = _T_116 | reset; // @[StrongEnum.scala 185:11]
  assign _T_119 = _T_118 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_120 = CastFromNonLit_25_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_122 = _T_120 | reset; // @[StrongEnum.scala 185:11]
  assign _T_123 = _T_122 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_124 = CastFromNonLit_26_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_126 = _T_124 | reset; // @[StrongEnum.scala 185:11]
  assign _T_127 = _T_126 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_128 = CastFromNonLit_27_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_130 = _T_128 | reset; // @[StrongEnum.scala 185:11]
  assign _T_131 = _T_130 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_132 = CastFromNonLit_28_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_134 = _T_132 | reset; // @[StrongEnum.scala 185:11]
  assign _T_135 = _T_134 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_136 = CastFromNonLit_29_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_138 = _T_136 | reset; // @[StrongEnum.scala 185:11]
  assign _T_139 = _T_138 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_140 = CastFromNonLit_30_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_142 = _T_140 | reset; // @[StrongEnum.scala 185:11]
  assign _T_143 = _T_142 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_144 = CastFromNonLit_31_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_146 = _T_144 | reset; // @[StrongEnum.scala 185:11]
  assign _T_147 = _T_146 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_148 = CastFromNonLit_32_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_150 = _T_148 | reset; // @[StrongEnum.scala 185:11]
  assign _T_151 = _T_150 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_152 = CastFromNonLit_33_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_154 = _T_152 | reset; // @[StrongEnum.scala 185:11]
  assign _T_155 = _T_154 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_156 = CastFromNonLit_34_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_158 = _T_156 | reset; // @[StrongEnum.scala 185:11]
  assign _T_159 = _T_158 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_160 = CastFromNonLit_35_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_162 = _T_160 | reset; // @[StrongEnum.scala 185:11]
  assign _T_163 = _T_162 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_164 = CastFromNonLit_36_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_166 = _T_164 | reset; // @[StrongEnum.scala 185:11]
  assign _T_167 = _T_166 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_168 = CastFromNonLit_37_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_170 = _T_168 | reset; // @[StrongEnum.scala 185:11]
  assign _T_171 = _T_170 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_172 = CastFromNonLit_38_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_174 = _T_172 | reset; // @[StrongEnum.scala 185:11]
  assign _T_175 = _T_174 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_176 = CastFromNonLit_39_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_178 = _T_176 | reset; // @[StrongEnum.scala 185:11]
  assign _T_179 = _T_178 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_180 = CastFromNonLit_40_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_182 = _T_180 | reset; // @[StrongEnum.scala 185:11]
  assign _T_183 = _T_182 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_184 = CastFromNonLit_41_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_186 = _T_184 | reset; // @[StrongEnum.scala 185:11]
  assign _T_187 = _T_186 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_188 = CastFromNonLit_42_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_190 = _T_188 | reset; // @[StrongEnum.scala 185:11]
  assign _T_191 = _T_190 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_192 = CastFromNonLit_43_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_194 = _T_192 | reset; // @[StrongEnum.scala 185:11]
  assign _T_195 = _T_194 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_196 = CastFromNonLit_44_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_198 = _T_196 | reset; // @[StrongEnum.scala 185:11]
  assign _T_199 = _T_198 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_200 = CastFromNonLit_45_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_202 = _T_200 | reset; // @[StrongEnum.scala 185:11]
  assign _T_203 = _T_202 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_204 = CastFromNonLit_46_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_206 = _T_204 | reset; // @[StrongEnum.scala 185:11]
  assign _T_207 = _T_206 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_208 = CastFromNonLit_47_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_210 = _T_208 | reset; // @[StrongEnum.scala 185:11]
  assign _T_211 = _T_210 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_212 = CastFromNonLit_48_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_214 = _T_212 | reset; // @[StrongEnum.scala 185:11]
  assign _T_215 = _T_214 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_216 = CastFromNonLit_49_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_218 = _T_216 | reset; // @[StrongEnum.scala 185:11]
  assign _T_219 = _T_218 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_220 = CastFromNonLit_50_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_222 = _T_220 | reset; // @[StrongEnum.scala 185:11]
  assign _T_223 = _T_222 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_224 = CastFromNonLit_51_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_226 = _T_224 | reset; // @[StrongEnum.scala 185:11]
  assign _T_227 = _T_226 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_228 = CastFromNonLit_52_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_230 = _T_228 | reset; // @[StrongEnum.scala 185:11]
  assign _T_231 = _T_230 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_232 = CastFromNonLit_53_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_234 = _T_232 | reset; // @[StrongEnum.scala 185:11]
  assign _T_235 = _T_234 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_236 = CastFromNonLit_54_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_238 = _T_236 | reset; // @[StrongEnum.scala 185:11]
  assign _T_239 = _T_238 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_240 = CastFromNonLit_55_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_242 = _T_240 | reset; // @[StrongEnum.scala 185:11]
  assign _T_243 = _T_242 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_244 = CastFromNonLit_56_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_246 = _T_244 | reset; // @[StrongEnum.scala 185:11]
  assign _T_247 = _T_246 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_248 = CastFromNonLit_57_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_250 = _T_248 | reset; // @[StrongEnum.scala 185:11]
  assign _T_251 = _T_250 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_252 = CastFromNonLit_58_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_254 = _T_252 | reset; // @[StrongEnum.scala 185:11]
  assign _T_255 = _T_254 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_256 = CastFromNonLit_59_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_258 = _T_256 | reset; // @[StrongEnum.scala 185:11]
  assign _T_259 = _T_258 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_260 = CastFromNonLit_60_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_262 = _T_260 | reset; // @[StrongEnum.scala 185:11]
  assign _T_263 = _T_262 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_264 = CastFromNonLit_61_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_266 = _T_264 | reset; // @[StrongEnum.scala 185:11]
  assign _T_267 = _T_266 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_268 = CastFromNonLit_62_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_270 = _T_268 | reset; // @[StrongEnum.scala 185:11]
  assign _T_271 = _T_270 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_272 = CastFromNonLit_63_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_274 = _T_272 | reset; // @[StrongEnum.scala 185:11]
  assign _T_275 = _T_274 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_276 = CastFromNonLit_64_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_278 = _T_276 | reset; // @[StrongEnum.scala 185:11]
  assign _T_279 = _T_278 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_280 = CastFromNonLit_65_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_282 = _T_280 | reset; // @[StrongEnum.scala 185:11]
  assign _T_283 = _T_282 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_284 = CastFromNonLit_66_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_286 = _T_284 | reset; // @[StrongEnum.scala 185:11]
  assign _T_287 = _T_286 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_288 = CastFromNonLit_67_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_290 = _T_288 | reset; // @[StrongEnum.scala 185:11]
  assign _T_291 = _T_290 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_292 = CastFromNonLit_68_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_294 = _T_292 | reset; // @[StrongEnum.scala 185:11]
  assign _T_295 = _T_294 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_296 = CastFromNonLit_69_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_298 = _T_296 | reset; // @[StrongEnum.scala 185:11]
  assign _T_299 = _T_298 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_300 = CastFromNonLit_70_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_302 = _T_300 | reset; // @[StrongEnum.scala 185:11]
  assign _T_303 = _T_302 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_304 = CastFromNonLit_71_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_306 = _T_304 | reset; // @[StrongEnum.scala 185:11]
  assign _T_307 = _T_306 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_308 = CastFromNonLit_72_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_310 = _T_308 | reset; // @[StrongEnum.scala 185:11]
  assign _T_311 = _T_310 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_312 = CastFromNonLit_73_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_314 = _T_312 | reset; // @[StrongEnum.scala 185:11]
  assign _T_315 = _T_314 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_316 = CastFromNonLit_74_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_318 = _T_316 | reset; // @[StrongEnum.scala 185:11]
  assign _T_319 = _T_318 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_320 = CastFromNonLit_75_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_322 = _T_320 | reset; // @[StrongEnum.scala 185:11]
  assign _T_323 = _T_322 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_324 = CastFromNonLit_76_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_326 = _T_324 | reset; // @[StrongEnum.scala 185:11]
  assign _T_327 = _T_326 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_328 = CastFromNonLit_77_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_330 = _T_328 | reset; // @[StrongEnum.scala 185:11]
  assign _T_331 = _T_330 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_332 = CastFromNonLit_78_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_334 = _T_332 | reset; // @[StrongEnum.scala 185:11]
  assign _T_335 = _T_334 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_336 = CastFromNonLit_79_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_338 = _T_336 | reset; // @[StrongEnum.scala 185:11]
  assign _T_339 = _T_338 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_340 = CastFromNonLit_80_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_342 = _T_340 | reset; // @[StrongEnum.scala 185:11]
  assign _T_343 = _T_342 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_344 = CastFromNonLit_81_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_346 = _T_344 | reset; // @[StrongEnum.scala 185:11]
  assign _T_347 = _T_346 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_348 = CastFromNonLit_82_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_350 = _T_348 | reset; // @[StrongEnum.scala 185:11]
  assign _T_351 = _T_350 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_352 = CastFromNonLit_83_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_354 = _T_352 | reset; // @[StrongEnum.scala 185:11]
  assign _T_355 = _T_354 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_356 = CastFromNonLit_84_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_358 = _T_356 | reset; // @[StrongEnum.scala 185:11]
  assign _T_359 = _T_358 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_360 = CastFromNonLit_85_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_362 = _T_360 | reset; // @[StrongEnum.scala 185:11]
  assign _T_363 = _T_362 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_364 = CastFromNonLit_86_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_366 = _T_364 | reset; // @[StrongEnum.scala 185:11]
  assign _T_367 = _T_366 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_368 = CastFromNonLit_87_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_370 = _T_368 | reset; // @[StrongEnum.scala 185:11]
  assign _T_371 = _T_370 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_372 = CastFromNonLit_88_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_374 = _T_372 | reset; // @[StrongEnum.scala 185:11]
  assign _T_375 = _T_374 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_376 = CastFromNonLit_89_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_378 = _T_376 | reset; // @[StrongEnum.scala 185:11]
  assign _T_379 = _T_378 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_380 = CastFromNonLit_90_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_382 = _T_380 | reset; // @[StrongEnum.scala 185:11]
  assign _T_383 = _T_382 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_384 = CastFromNonLit_91_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_386 = _T_384 | reset; // @[StrongEnum.scala 185:11]
  assign _T_387 = _T_386 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_388 = CastFromNonLit_92_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_390 = _T_388 | reset; // @[StrongEnum.scala 185:11]
  assign _T_391 = _T_390 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_392 = CastFromNonLit_93_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_394 = _T_392 | reset; // @[StrongEnum.scala 185:11]
  assign _T_395 = _T_394 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_396 = CastFromNonLit_94_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_398 = _T_396 | reset; // @[StrongEnum.scala 185:11]
  assign _T_399 = _T_398 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_400 = CastFromNonLit_95_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_402 = _T_400 | reset; // @[StrongEnum.scala 185:11]
  assign _T_403 = _T_402 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_404 = CastFromNonLit_96_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_406 = _T_404 | reset; // @[StrongEnum.scala 185:11]
  assign _T_407 = _T_406 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_408 = CastFromNonLit_97_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_410 = _T_408 | reset; // @[StrongEnum.scala 185:11]
  assign _T_411 = _T_410 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_412 = CastFromNonLit_98_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_414 = _T_412 | reset; // @[StrongEnum.scala 185:11]
  assign _T_415 = _T_414 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_416 = CastFromNonLit_99_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_418 = _T_416 | reset; // @[StrongEnum.scala 185:11]
  assign _T_419 = _T_418 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_420 = CastFromNonLit_100_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_422 = _T_420 | reset; // @[StrongEnum.scala 185:11]
  assign _T_423 = _T_422 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_424 = CastFromNonLit_101_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_426 = _T_424 | reset; // @[StrongEnum.scala 185:11]
  assign _T_427 = _T_426 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_428 = CastFromNonLit_102_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_430 = _T_428 | reset; // @[StrongEnum.scala 185:11]
  assign _T_431 = _T_430 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_432 = CastFromNonLit_103_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_434 = _T_432 | reset; // @[StrongEnum.scala 185:11]
  assign _T_435 = _T_434 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_436 = CastFromNonLit_104_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_438 = _T_436 | reset; // @[StrongEnum.scala 185:11]
  assign _T_439 = _T_438 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_440 = CastFromNonLit_105_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_442 = _T_440 | reset; // @[StrongEnum.scala 185:11]
  assign _T_443 = _T_442 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_444 = CastFromNonLit_106_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_446 = _T_444 | reset; // @[StrongEnum.scala 185:11]
  assign _T_447 = _T_446 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_448 = CastFromNonLit_107_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_450 = _T_448 | reset; // @[StrongEnum.scala 185:11]
  assign _T_451 = _T_450 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_452 = CastFromNonLit_108_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_454 = _T_452 | reset; // @[StrongEnum.scala 185:11]
  assign _T_455 = _T_454 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_456 = CastFromNonLit_109_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_458 = _T_456 | reset; // @[StrongEnum.scala 185:11]
  assign _T_459 = _T_458 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_460 = CastFromNonLit_110_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_462 = _T_460 | reset; // @[StrongEnum.scala 185:11]
  assign _T_463 = _T_462 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_464 = CastFromNonLit_111_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_466 = _T_464 | reset; // @[StrongEnum.scala 185:11]
  assign _T_467 = _T_466 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_468 = CastFromNonLit_112_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_470 = _T_468 | reset; // @[StrongEnum.scala 185:11]
  assign _T_471 = _T_470 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_472 = CastFromNonLit_113_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_474 = _T_472 | reset; // @[StrongEnum.scala 185:11]
  assign _T_475 = _T_474 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_476 = CastFromNonLit_114_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_478 = _T_476 | reset; // @[StrongEnum.scala 185:11]
  assign _T_479 = _T_478 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_480 = CastFromNonLit_115_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_482 = _T_480 | reset; // @[StrongEnum.scala 185:11]
  assign _T_483 = _T_482 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_484 = CastFromNonLit_116_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_486 = _T_484 | reset; // @[StrongEnum.scala 185:11]
  assign _T_487 = _T_486 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_488 = CastFromNonLit_117_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_490 = _T_488 | reset; // @[StrongEnum.scala 185:11]
  assign _T_491 = _T_490 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_492 = CastFromNonLit_118_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_494 = _T_492 | reset; // @[StrongEnum.scala 185:11]
  assign _T_495 = _T_494 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_496 = CastFromNonLit_119_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_498 = _T_496 | reset; // @[StrongEnum.scala 185:11]
  assign _T_499 = _T_498 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_500 = CastFromNonLit_120_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_502 = _T_500 | reset; // @[StrongEnum.scala 185:11]
  assign _T_503 = _T_502 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_504 = CastFromNonLit_121_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_506 = _T_504 | reset; // @[StrongEnum.scala 185:11]
  assign _T_507 = _T_506 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_508 = CastFromNonLit_122_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_510 = _T_508 | reset; // @[StrongEnum.scala 185:11]
  assign _T_511 = _T_510 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_512 = CastFromNonLit_123_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_514 = _T_512 | reset; // @[StrongEnum.scala 185:11]
  assign _T_515 = _T_514 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_516 = CastFromNonLit_124_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_518 = _T_516 | reset; // @[StrongEnum.scala 185:11]
  assign _T_519 = _T_518 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_520 = CastFromNonLit_125_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_522 = _T_520 | reset; // @[StrongEnum.scala 185:11]
  assign _T_523 = _T_522 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_524 = CastFromNonLit_126_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_526 = _T_524 | reset; // @[StrongEnum.scala 185:11]
  assign _T_527 = _T_526 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_528 = CastFromNonLit_127_io_valid == 1'h0; // @[StrongEnum.scala 185:25]
  assign _T_530 = _T_528 | reset; // @[StrongEnum.scala 185:11]
  assign _T_531 = _T_530 == 1'h0; // @[StrongEnum.scala 185:11]
  assign _T_533 = reset == 1'h0; // @[StrongEnum.scala 188:7]
  assign CastFromNonLit_io_in = 7'h0; // @[StrongEnum.scala 172:15]
  assign CastFromNonLit_1_io_in = 7'h1; // @[StrongEnum.scala 172:15]
  assign CastFromNonLit_2_io_in = 7'h2; // @[StrongEnum.scala 172:15]
  assign CastFromNonLit_3_io_in = 7'h64; // @[StrongEnum.scala 172:15]
  assign CastFromNonLit_4_io_in = 7'h65; // @[StrongEnum.scala 172:15]
  assign CastFromNonLit_5_io_in = 7'h3; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_6_io_in = 7'h4; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_7_io_in = 7'h5; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_8_io_in = 7'h6; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_9_io_in = 7'h7; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_10_io_in = 7'h8; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_11_io_in = 7'h9; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_12_io_in = 7'ha; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_13_io_in = 7'hb; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_14_io_in = 7'hc; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_15_io_in = 7'hd; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_16_io_in = 7'he; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_17_io_in = 7'hf; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_18_io_in = 7'h10; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_19_io_in = 7'h11; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_20_io_in = 7'h12; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_21_io_in = 7'h13; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_22_io_in = 7'h14; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_23_io_in = 7'h15; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_24_io_in = 7'h16; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_25_io_in = 7'h17; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_26_io_in = 7'h18; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_27_io_in = 7'h19; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_28_io_in = 7'h1a; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_29_io_in = 7'h1b; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_30_io_in = 7'h1c; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_31_io_in = 7'h1d; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_32_io_in = 7'h1e; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_33_io_in = 7'h1f; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_34_io_in = 7'h20; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_35_io_in = 7'h21; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_36_io_in = 7'h22; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_37_io_in = 7'h23; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_38_io_in = 7'h24; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_39_io_in = 7'h25; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_40_io_in = 7'h26; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_41_io_in = 7'h27; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_42_io_in = 7'h28; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_43_io_in = 7'h29; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_44_io_in = 7'h2a; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_45_io_in = 7'h2b; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_46_io_in = 7'h2c; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_47_io_in = 7'h2d; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_48_io_in = 7'h2e; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_49_io_in = 7'h2f; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_50_io_in = 7'h30; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_51_io_in = 7'h31; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_52_io_in = 7'h32; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_53_io_in = 7'h33; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_54_io_in = 7'h34; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_55_io_in = 7'h35; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_56_io_in = 7'h36; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_57_io_in = 7'h37; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_58_io_in = 7'h38; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_59_io_in = 7'h39; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_60_io_in = 7'h3a; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_61_io_in = 7'h3b; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_62_io_in = 7'h3c; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_63_io_in = 7'h3d; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_64_io_in = 7'h3e; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_65_io_in = 7'h3f; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_66_io_in = 7'h40; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_67_io_in = 7'h41; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_68_io_in = 7'h42; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_69_io_in = 7'h43; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_70_io_in = 7'h44; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_71_io_in = 7'h45; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_72_io_in = 7'h46; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_73_io_in = 7'h47; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_74_io_in = 7'h48; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_75_io_in = 7'h49; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_76_io_in = 7'h4a; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_77_io_in = 7'h4b; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_78_io_in = 7'h4c; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_79_io_in = 7'h4d; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_80_io_in = 7'h4e; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_81_io_in = 7'h4f; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_82_io_in = 7'h50; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_83_io_in = 7'h51; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_84_io_in = 7'h52; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_85_io_in = 7'h53; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_86_io_in = 7'h54; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_87_io_in = 7'h55; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_88_io_in = 7'h56; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_89_io_in = 7'h57; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_90_io_in = 7'h58; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_91_io_in = 7'h59; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_92_io_in = 7'h5a; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_93_io_in = 7'h5b; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_94_io_in = 7'h5c; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_95_io_in = 7'h5d; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_96_io_in = 7'h5e; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_97_io_in = 7'h5f; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_98_io_in = 7'h60; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_99_io_in = 7'h61; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_100_io_in = 7'h62; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_101_io_in = 7'h63; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_102_io_in = 7'h66; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_103_io_in = 7'h67; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_104_io_in = 7'h68; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_105_io_in = 7'h69; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_106_io_in = 7'h6a; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_107_io_in = 7'h6b; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_108_io_in = 7'h6c; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_109_io_in = 7'h6d; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_110_io_in = 7'h6e; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_111_io_in = 7'h6f; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_112_io_in = 7'h70; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_113_io_in = 7'h71; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_114_io_in = 7'h72; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_115_io_in = 7'h73; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_116_io_in = 7'h74; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_117_io_in = 7'h75; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_118_io_in = 7'h76; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_119_io_in = 7'h77; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_120_io_in = 7'h78; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_121_io_in = 7'h79; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_122_io_in = 7'h7a; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_123_io_in = 7'h7b; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_124_io_in = 7'h7c; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_125_io_in = 7'h7d; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_126_io_in = 7'h7e; // @[StrongEnum.scala 183:15]
  assign CastFromNonLit_127_io_in = 7'h7f; // @[StrongEnum.scala 183:15]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:173 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 173:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3) begin
          $fatal; // @[StrongEnum.scala 173:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:174 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 174:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7) begin
          $fatal; // @[StrongEnum.scala 174:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:173 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 173:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_11) begin
          $fatal; // @[StrongEnum.scala 173:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:174 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 174:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_15) begin
          $fatal; // @[StrongEnum.scala 174:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:173 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 173:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_19) begin
          $fatal; // @[StrongEnum.scala 173:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_23) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:174 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 174:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_23) begin
          $fatal; // @[StrongEnum.scala 174:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_27) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:173 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 173:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_27) begin
          $fatal; // @[StrongEnum.scala 173:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_31) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:174 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 174:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_31) begin
          $fatal; // @[StrongEnum.scala 174:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:173 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 173:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_35) begin
          $fatal; // @[StrongEnum.scala 173:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:174 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 174:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_39) begin
          $fatal; // @[StrongEnum.scala 174:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_43) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_43) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_47) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_47) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_51) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_51) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_55) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_55) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_59) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_59) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_63) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_67) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_67) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_71) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_71) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_75) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_75) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_79) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_79) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_83) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_83) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_87) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_87) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_91) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_91) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_95) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_95) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_99) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_99) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_103) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_103) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_107) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_107) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_111) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_111) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_115) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_115) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_119) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_119) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_123) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_123) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_127) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_127) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_131) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_135) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_135) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_139) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_139) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_143) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_143) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_147) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_147) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_151) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_151) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_155) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_155) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_159) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_159) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_163) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_163) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_167) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_167) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_171) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_171) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_175) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_175) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_179) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_179) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_183) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_183) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_187) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_187) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_191) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_191) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_195) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_195) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_199) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_199) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_203) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_203) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_207) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_207) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_211) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_211) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_215) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_215) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_219) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_223) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_223) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_227) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_227) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_231) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_231) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_235) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_235) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_239) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_239) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_243) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_243) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_247) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_247) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_251) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_251) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_255) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_255) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_259) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_259) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_263) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_263) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_267) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_267) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_271) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_271) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_275) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_275) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_279) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_279) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_283) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_283) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_287) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_287) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_291) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_291) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_295) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_295) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_299) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_299) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_303) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_303) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_307) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_307) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_311) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_311) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_315) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_315) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_319) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_319) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_323) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_323) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_327) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_327) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_331) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_331) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_335) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_335) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_339) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_339) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_343) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_343) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_347) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_347) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_351) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_351) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_355) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_355) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_359) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_359) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_363) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_363) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_367) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_367) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_371) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_371) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_375) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_375) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_379) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_379) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_383) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_383) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_387) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_387) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_391) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_391) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_395) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_395) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_399) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_399) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_403) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_403) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_407) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_407) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_411) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_411) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_415) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_415) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_419) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_419) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_423) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_423) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_427) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_427) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_431) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_431) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_435) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_435) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_439) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_439) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_443) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_443) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_447) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_447) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_451) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_451) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_455) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_455) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_459) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_459) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_463) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_463) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_467) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_467) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_471) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_471) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_475) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_475) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_479) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_479) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_483) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_483) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_487) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_487) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_491) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_491) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_495) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_495) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_499) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_499) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_503) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_503) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_507) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_507) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_511) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_511) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_515) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_515) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_519) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_519) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_523) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_523) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_527) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_527) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_531) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:185 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 185:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_531) begin
          $fatal; // @[StrongEnum.scala 185:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_533) begin
          $finish; // @[StrongEnum.scala 188:7]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
