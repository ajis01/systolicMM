module RoundAnyRawFNToRecFN(
  input         io_in_isZero,
  input  [7:0]  io_in_sExp,
  input  [32:0] io_in_sig,
  output [64:0] io_out
);
  wire [11:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] _T_3; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire [55:0] adjustedSig; // @[RoundAnyRawFNToRecFN.scala 112:22]
  wire [12:0] _T_6; // @[RoundAnyRawFNToRecFN.scala 134:55]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 134:55]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 138:28]
  wire [11:0] _T_22; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [12:0] _T_48; // @[Cat.scala 29:58]
  assign _GEN_0 = {{4{io_in_sExp[7]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign _T_3 = $signed(_GEN_0) + 12'sh7c0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_T_3[11:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign adjustedSig = {io_in_sig, 23'h0}; // @[RoundAnyRawFNToRecFN.scala 112:22]
  assign _T_6 = {{1'd0}, sAdjustedExp[11:0]}; // @[RoundAnyRawFNToRecFN.scala 134:55]
  assign common_expOut = _T_6[11:0]; // @[RoundAnyRawFNToRecFN.scala 134:55]
  assign common_fractOut = adjustedSig[53:2]; // @[RoundAnyRawFNToRecFN.scala 138:28]
  assign _T_22 = io_in_isZero ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign expOut = common_expOut & ~_T_22; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign fractOut = io_in_isZero ? 52'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _T_48 = {1'h0,expOut}; // @[Cat.scala 29:58]
  assign io_out = {_T_48,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
endmodule
module INToRecFN(
  input  [31:0] io_in,
  output [64:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire [7:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [32:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [63:0] _T_5; // @[Cat.scala 29:58]
  wire [4:0] _T_39; // @[Mux.scala 47:69]
  wire [4:0] _T_40; // @[Mux.scala 47:69]
  wire [4:0] _T_41; // @[Mux.scala 47:69]
  wire [4:0] _T_42; // @[Mux.scala 47:69]
  wire [4:0] _T_43; // @[Mux.scala 47:69]
  wire [4:0] _T_44; // @[Mux.scala 47:69]
  wire [4:0] _T_45; // @[Mux.scala 47:69]
  wire [4:0] _T_46; // @[Mux.scala 47:69]
  wire [4:0] _T_47; // @[Mux.scala 47:69]
  wire [4:0] _T_48; // @[Mux.scala 47:69]
  wire [4:0] _T_49; // @[Mux.scala 47:69]
  wire [4:0] _T_50; // @[Mux.scala 47:69]
  wire [4:0] _T_51; // @[Mux.scala 47:69]
  wire [4:0] _T_52; // @[Mux.scala 47:69]
  wire [4:0] _T_53; // @[Mux.scala 47:69]
  wire [4:0] _T_54; // @[Mux.scala 47:69]
  wire [4:0] _T_55; // @[Mux.scala 47:69]
  wire [4:0] _T_56; // @[Mux.scala 47:69]
  wire [4:0] _T_57; // @[Mux.scala 47:69]
  wire [4:0] _T_58; // @[Mux.scala 47:69]
  wire [4:0] _T_59; // @[Mux.scala 47:69]
  wire [4:0] _T_60; // @[Mux.scala 47:69]
  wire [4:0] _T_61; // @[Mux.scala 47:69]
  wire [4:0] _T_62; // @[Mux.scala 47:69]
  wire [4:0] _T_63; // @[Mux.scala 47:69]
  wire [4:0] _T_64; // @[Mux.scala 47:69]
  wire [4:0] _T_65; // @[Mux.scala 47:69]
  wire [4:0] _T_66; // @[Mux.scala 47:69]
  wire [4:0] _T_67; // @[Mux.scala 47:69]
  wire [4:0] _T_68; // @[Mux.scala 47:69]
  wire [4:0] _T_69; // @[Mux.scala 47:69]
  wire [62:0] _GEN_0; // @[rawFloatFromIN.scala 55:22]
  wire [62:0] _T_70; // @[rawFloatFromIN.scala 55:22]
  wire [6:0] _T_76; // @[Cat.scala 29:58]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign _T_5 = {32'h0,io_in}; // @[Cat.scala 29:58]
  assign _T_39 = _T_5[1] ? 5'h1e : 5'h1f; // @[Mux.scala 47:69]
  assign _T_40 = _T_5[2] ? 5'h1d : _T_39; // @[Mux.scala 47:69]
  assign _T_41 = _T_5[3] ? 5'h1c : _T_40; // @[Mux.scala 47:69]
  assign _T_42 = _T_5[4] ? 5'h1b : _T_41; // @[Mux.scala 47:69]
  assign _T_43 = _T_5[5] ? 5'h1a : _T_42; // @[Mux.scala 47:69]
  assign _T_44 = _T_5[6] ? 5'h19 : _T_43; // @[Mux.scala 47:69]
  assign _T_45 = _T_5[7] ? 5'h18 : _T_44; // @[Mux.scala 47:69]
  assign _T_46 = _T_5[8] ? 5'h17 : _T_45; // @[Mux.scala 47:69]
  assign _T_47 = _T_5[9] ? 5'h16 : _T_46; // @[Mux.scala 47:69]
  assign _T_48 = _T_5[10] ? 5'h15 : _T_47; // @[Mux.scala 47:69]
  assign _T_49 = _T_5[11] ? 5'h14 : _T_48; // @[Mux.scala 47:69]
  assign _T_50 = _T_5[12] ? 5'h13 : _T_49; // @[Mux.scala 47:69]
  assign _T_51 = _T_5[13] ? 5'h12 : _T_50; // @[Mux.scala 47:69]
  assign _T_52 = _T_5[14] ? 5'h11 : _T_51; // @[Mux.scala 47:69]
  assign _T_53 = _T_5[15] ? 5'h10 : _T_52; // @[Mux.scala 47:69]
  assign _T_54 = _T_5[16] ? 5'hf : _T_53; // @[Mux.scala 47:69]
  assign _T_55 = _T_5[17] ? 5'he : _T_54; // @[Mux.scala 47:69]
  assign _T_56 = _T_5[18] ? 5'hd : _T_55; // @[Mux.scala 47:69]
  assign _T_57 = _T_5[19] ? 5'hc : _T_56; // @[Mux.scala 47:69]
  assign _T_58 = _T_5[20] ? 5'hb : _T_57; // @[Mux.scala 47:69]
  assign _T_59 = _T_5[21] ? 5'ha : _T_58; // @[Mux.scala 47:69]
  assign _T_60 = _T_5[22] ? 5'h9 : _T_59; // @[Mux.scala 47:69]
  assign _T_61 = _T_5[23] ? 5'h8 : _T_60; // @[Mux.scala 47:69]
  assign _T_62 = _T_5[24] ? 5'h7 : _T_61; // @[Mux.scala 47:69]
  assign _T_63 = _T_5[25] ? 5'h6 : _T_62; // @[Mux.scala 47:69]
  assign _T_64 = _T_5[26] ? 5'h5 : _T_63; // @[Mux.scala 47:69]
  assign _T_65 = _T_5[27] ? 5'h4 : _T_64; // @[Mux.scala 47:69]
  assign _T_66 = _T_5[28] ? 5'h3 : _T_65; // @[Mux.scala 47:69]
  assign _T_67 = _T_5[29] ? 5'h2 : _T_66; // @[Mux.scala 47:69]
  assign _T_68 = _T_5[30] ? 5'h1 : _T_67; // @[Mux.scala 47:69]
  assign _T_69 = _T_5[31] ? 5'h0 : _T_68; // @[Mux.scala 47:69]
  assign _GEN_0 = {{31'd0}, _T_5[31:0]}; // @[rawFloatFromIN.scala 55:22]
  assign _T_70 = _GEN_0 << _T_69; // @[rawFloatFromIN.scala 55:22]
  assign _T_76 = {2'h2,~_T_69}; // @[Cat.scala 29:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_70[31]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_76)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_70[31:0]}; // @[INToRecFN.scala 69:44]
endmodule
module ValExec_UI32ToRecF64(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  input  [63:0] io_expected_out,
  input  [4:0]  io_expected_exceptionFlags,
  output [64:0] io_expected_recOut,
  output [64:0] io_actual_out,
  output [4:0]  io_actual_exceptionFlags,
  output        io_check,
  output        io_pass
);
  wire [31:0] iNToRecFN_io_in; // @[ValExec_INToRecFN.scala 66:27]
  wire [64:0] iNToRecFN_io_out; // @[ValExec_INToRecFN.scala 66:27]
  wire  _T_3; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_57; // @[Mux.scala 47:69]
  wire [5:0] _T_58; // @[Mux.scala 47:69]
  wire [5:0] _T_59; // @[Mux.scala 47:69]
  wire [5:0] _T_60; // @[Mux.scala 47:69]
  wire [5:0] _T_61; // @[Mux.scala 47:69]
  wire [5:0] _T_62; // @[Mux.scala 47:69]
  wire [5:0] _T_63; // @[Mux.scala 47:69]
  wire [5:0] _T_64; // @[Mux.scala 47:69]
  wire [5:0] _T_65; // @[Mux.scala 47:69]
  wire [5:0] _T_66; // @[Mux.scala 47:69]
  wire [5:0] _T_67; // @[Mux.scala 47:69]
  wire [5:0] _T_68; // @[Mux.scala 47:69]
  wire [5:0] _T_69; // @[Mux.scala 47:69]
  wire [5:0] _T_70; // @[Mux.scala 47:69]
  wire [5:0] _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_107; // @[Mux.scala 47:69]
  wire [114:0] _GEN_0; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_108; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_110; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_1; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_111; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_112; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_113; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_114; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_116; // @[rawFloatFromFN.scala 59:15]
  wire  _T_117; // @[rawFloatFromFN.scala 62:34]
  wire  _T_119; // @[rawFloatFromFN.scala 63:62]
  wire  _T_122; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_125; // @[rawFloatFromFN.scala 70:48]
  wire [51:0] _T_127; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_129; // @[Cat.scala 29:58]
  wire [2:0] _T_131; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_133; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_136; // @[Cat.scala 29:58]
  wire [3:0] _T_137; // @[Cat.scala 29:58]
  wire  _T_142; // @[tests.scala 48:26]
  wire  _T_144; // @[tests.scala 48:55]
  wire  _T_145; // @[tests.scala 48:39]
  wire  _T_146; // @[tests.scala 49:20]
  wire  _T_149; // @[tests.scala 49:54]
  wire  _T_150; // @[tests.scala 49:31]
  wire  _T_152; // @[tests.scala 50:30]
  wire  _T_154; // @[tests.scala 50:66]
  wire  _T_155; // @[tests.scala 50:16]
  wire  _T_156; // @[tests.scala 48:12]
  wire  _T_157; // @[ValExec_INToRecFN.scala 80:35]
  INToRecFN iNToRecFN ( // @[ValExec_INToRecFN.scala 66:27]
    .io_in(iNToRecFN_io_in),
    .io_out(iNToRecFN_io_out)
  );
  assign _T_3 = io_expected_out[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign _T_4 = io_expected_out[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _T_57 = io_expected_out[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _T_58 = io_expected_out[2] ? 6'h31 : _T_57; // @[Mux.scala 47:69]
  assign _T_59 = io_expected_out[3] ? 6'h30 : _T_58; // @[Mux.scala 47:69]
  assign _T_60 = io_expected_out[4] ? 6'h2f : _T_59; // @[Mux.scala 47:69]
  assign _T_61 = io_expected_out[5] ? 6'h2e : _T_60; // @[Mux.scala 47:69]
  assign _T_62 = io_expected_out[6] ? 6'h2d : _T_61; // @[Mux.scala 47:69]
  assign _T_63 = io_expected_out[7] ? 6'h2c : _T_62; // @[Mux.scala 47:69]
  assign _T_64 = io_expected_out[8] ? 6'h2b : _T_63; // @[Mux.scala 47:69]
  assign _T_65 = io_expected_out[9] ? 6'h2a : _T_64; // @[Mux.scala 47:69]
  assign _T_66 = io_expected_out[10] ? 6'h29 : _T_65; // @[Mux.scala 47:69]
  assign _T_67 = io_expected_out[11] ? 6'h28 : _T_66; // @[Mux.scala 47:69]
  assign _T_68 = io_expected_out[12] ? 6'h27 : _T_67; // @[Mux.scala 47:69]
  assign _T_69 = io_expected_out[13] ? 6'h26 : _T_68; // @[Mux.scala 47:69]
  assign _T_70 = io_expected_out[14] ? 6'h25 : _T_69; // @[Mux.scala 47:69]
  assign _T_71 = io_expected_out[15] ? 6'h24 : _T_70; // @[Mux.scala 47:69]
  assign _T_72 = io_expected_out[16] ? 6'h23 : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = io_expected_out[17] ? 6'h22 : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = io_expected_out[18] ? 6'h21 : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = io_expected_out[19] ? 6'h20 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = io_expected_out[20] ? 6'h1f : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = io_expected_out[21] ? 6'h1e : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = io_expected_out[22] ? 6'h1d : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = io_expected_out[23] ? 6'h1c : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = io_expected_out[24] ? 6'h1b : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = io_expected_out[25] ? 6'h1a : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = io_expected_out[26] ? 6'h19 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = io_expected_out[27] ? 6'h18 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = io_expected_out[28] ? 6'h17 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = io_expected_out[29] ? 6'h16 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = io_expected_out[30] ? 6'h15 : _T_85; // @[Mux.scala 47:69]
  assign _T_87 = io_expected_out[31] ? 6'h14 : _T_86; // @[Mux.scala 47:69]
  assign _T_88 = io_expected_out[32] ? 6'h13 : _T_87; // @[Mux.scala 47:69]
  assign _T_89 = io_expected_out[33] ? 6'h12 : _T_88; // @[Mux.scala 47:69]
  assign _T_90 = io_expected_out[34] ? 6'h11 : _T_89; // @[Mux.scala 47:69]
  assign _T_91 = io_expected_out[35] ? 6'h10 : _T_90; // @[Mux.scala 47:69]
  assign _T_92 = io_expected_out[36] ? 6'hf : _T_91; // @[Mux.scala 47:69]
  assign _T_93 = io_expected_out[37] ? 6'he : _T_92; // @[Mux.scala 47:69]
  assign _T_94 = io_expected_out[38] ? 6'hd : _T_93; // @[Mux.scala 47:69]
  assign _T_95 = io_expected_out[39] ? 6'hc : _T_94; // @[Mux.scala 47:69]
  assign _T_96 = io_expected_out[40] ? 6'hb : _T_95; // @[Mux.scala 47:69]
  assign _T_97 = io_expected_out[41] ? 6'ha : _T_96; // @[Mux.scala 47:69]
  assign _T_98 = io_expected_out[42] ? 6'h9 : _T_97; // @[Mux.scala 47:69]
  assign _T_99 = io_expected_out[43] ? 6'h8 : _T_98; // @[Mux.scala 47:69]
  assign _T_100 = io_expected_out[44] ? 6'h7 : _T_99; // @[Mux.scala 47:69]
  assign _T_101 = io_expected_out[45] ? 6'h6 : _T_100; // @[Mux.scala 47:69]
  assign _T_102 = io_expected_out[46] ? 6'h5 : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = io_expected_out[47] ? 6'h4 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = io_expected_out[48] ? 6'h3 : _T_103; // @[Mux.scala 47:69]
  assign _T_105 = io_expected_out[49] ? 6'h2 : _T_104; // @[Mux.scala 47:69]
  assign _T_106 = io_expected_out[50] ? 6'h1 : _T_105; // @[Mux.scala 47:69]
  assign _T_107 = io_expected_out[51] ? 6'h0 : _T_106; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, io_expected_out[51:0]}; // @[rawFloatFromFN.scala 54:36]
  assign _T_108 = _GEN_0 << _T_107; // @[rawFloatFromFN.scala 54:36]
  assign _T_110 = {_T_108[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_1 = {{6'd0}, _T_107}; // @[rawFloatFromFN.scala 57:26]
  assign _T_111 = _GEN_1 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _T_112 = _T_3 ? _T_111 : {{1'd0}, io_expected_out[62:52]}; // @[rawFloatFromFN.scala 56:16]
  assign _T_113 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_2 = {{9'd0}, _T_113}; // @[rawFloatFromFN.scala 60:22]
  assign _T_114 = 11'h400 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_3 = {{1'd0}, _T_114}; // @[rawFloatFromFN.scala 59:15]
  assign _T_116 = _T_112 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  assign _T_117 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  assign _T_119 = _T_116[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign _T_122 = _T_119 & ~_T_4; // @[rawFloatFromFN.scala 66:33]
  assign _T_125 = {1'b0,$signed(_T_116)}; // @[rawFloatFromFN.scala 70:48]
  assign _T_127 = _T_3 ? _T_110 : io_expected_out[51:0]; // @[rawFloatFromFN.scala 72:42]
  assign _T_129 = {1'h0,~_T_117,_T_127}; // @[Cat.scala 29:58]
  assign _T_131 = _T_117 ? 3'h0 : _T_125[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_4 = {{2'd0}, _T_122}; // @[recFNFromFN.scala 48:79]
  assign _T_133 = _T_131 | _GEN_4; // @[recFNFromFN.scala 48:79]
  assign _T_136 = {_T_125[8:0],_T_129[51:0]}; // @[Cat.scala 29:58]
  assign _T_137 = {io_expected_out[63],_T_133}; // @[Cat.scala 29:58]
  assign _T_142 = io_actual_out[63:61] == 3'h0; // @[tests.scala 48:26]
  assign _T_144 = io_actual_out[63:61] == 3'h7; // @[tests.scala 48:55]
  assign _T_145 = _T_142 | _T_144; // @[tests.scala 48:39]
  assign _T_146 = io_actual_out[64:61] == io_expected_recOut[64:61]; // @[tests.scala 49:20]
  assign _T_149 = io_actual_out[51:0] == io_expected_recOut[51:0]; // @[tests.scala 49:54]
  assign _T_150 = _T_146 & _T_149; // @[tests.scala 49:31]
  assign _T_152 = io_actual_out[63:61] == 3'h6; // @[tests.scala 50:30]
  assign _T_154 = io_actual_out == io_expected_recOut; // @[tests.scala 50:66]
  assign _T_155 = _T_152 ? _T_146 : _T_154; // @[tests.scala 50:16]
  assign _T_156 = _T_145 ? _T_150 : _T_155; // @[tests.scala 48:12]
  assign _T_157 = io_actual_exceptionFlags == io_expected_exceptionFlags; // @[ValExec_INToRecFN.scala 80:35]
  assign io_expected_recOut = {_T_137,_T_136}; // @[ValExec_INToRecFN.scala 72:24]
  assign io_actual_out = iNToRecFN_io_out; // @[ValExec_INToRecFN.scala 74:19]
  assign io_actual_exceptionFlags = 5'h0; // @[ValExec_INToRecFN.scala 75:30]
  assign io_check = 1'h1; // @[ValExec_INToRecFN.scala 77:14]
  assign io_pass = _T_156 & _T_157; // @[ValExec_INToRecFN.scala 78:13]
  assign iNToRecFN_io_in = io_in; // @[ValExec_INToRecFN.scala 68:21]
endmodule
