module SinglePrintfTester(
  input   clock,
  input   reset
);
  wire  _T_1; // @[Printf.scala 10:9]
  assign _T_1 = reset == 1'h0; // @[Printf.scala 10:9]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"x=%x",8'hfe); // @[Printf.scala 10:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1) begin
          $finish; // @[Printf.scala 11:7]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
